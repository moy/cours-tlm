XlxV37EB    14ee     61exڽXko9�ί�J"m�
�C*i*���Hi��j����1`�`��V���\�!��]�Ηƾ����*��^�J��q�\��VD������3֚��x��T���V{��^qrB����׍�r^8'���cJ���5[�U����:&a���2򙕥\��wwM�&�X5����z������Q�Γ��GV:i�2���U���U��*G^>z���BiG�5�U�;)�۾�%����)�7v$�2�L��2�X9oU/�2f*��e:��I�$��-a��3GbB=I��qy^dR��!��XV&J���dBif]&�'o�%x�#�6
�D�s%��J9e��L�V{w��;=2����d6�` ��A&,l�X��i"��dZߔ���3熭�\� "�����؋r}(�ߤd#����RgYG���Ӟp���9�ڬ�G/Q�i��F��f����"M���_鏩���}��WtO���P�0��T:J2�]ɟ�#�E�ɱL���Y�f�"�Qj���u.�.��L$ץD�<N����x/gϥ�yί�K릵�E"��3�beQ�T^6(�J�҄}9#G��rFZg�y��x����f�@��Q��K��̱��fDB3����l�+�]��8��ǋ�&u�E)�D��%ݎ��H9�#�ϙWx���Q4k���Y��DTXeP&Z����s|]}���Z�I��H����o���s�>�T"���L�u��t��(]dU�a��;�^��+¯ҙ&>����}�Vt���`�X��f�v��y��6��&��ȱrs�p,���{Ff7���oV��S�|F
;i䦇�(Tjo+/k��IYd��<M���K1�n�4z��*Uc��P�@NP�]ce��w��\
�V��f�\*J�D��[7V�������"xX�?� 7貐H-��6�����qAC&�F���OR������VAmӣ|	|x�\k.H�Ucgn�\�Y˳叢���r���LJ<��'��̨ ��T&�>��V���cv���ҁ���|�wi�4,P��imfEe�<ŧ�PhW^��Sh9�8-F��������zHaO�`n�\!s0:����ֻ4�6¨T@��
�j\�\5[�βkS�9`�2���}*��uy۾��ow�������~�"Q=�oEj�Z���#<U������[��yUE�-,�l���Ŧ|�$�o�U�Ci	�`��tXb�:�oIB�gA�8�z-,��roM7���h�C��=�=��T�h�z%���%���˧��t3<�f��@FL���F�������<:ܔ����r>7�]��y��V��#a�Ѧ�aw)OB0?U�(�a7�;�{�k�q��z��`4�5���\L�'��@A},���a;����QC��N��/wߚ�݋n����"�Qy�i ���Mg�Pyu�W菥��Q��� ������`V� b�ܨ���;�J����⪠�m�R�~�O����M��poޯg�]�s���`�zP���4��r��!�B�<� ���4�