XlxV37EB    fa00    28c7x��=ks�8���+pޫ�=��%;�l��*Y��Z�O��ٚb�l�"��r���A`%���.f���n ���7o&����O�i�l����!�п�O�>����"��}���~@��Q������#�=��9�t�ey�eQ�#�q���%�3�]9�]Ao^�q��.Jgwq�g�:�/�&m�����'��4����/�"^>�F�r��z�bJq��<˾lҥ���x���=�$���
��Y�,K��y{p�O�fi��������k<��9Z��gY��Y�b�=��������7�
�%����M�O����/х�:�K�J��6I�%��%��$}����~Ft�v��9�@aO�4�ŀp�<�0pGo:]
�c��'���ߦ�z/o��|��,��G9A�a=���!�^gF�V�dP���F�x��x��N�<�8������h9_���0������U0�2�Tv4����w�ŷ�h�}BП���n�5[$�ov�5[|�}���ㇿ����q��oT�.��P��/�������$42v)��xI�(Za3��_/|	�l
9F�Q�K���1�?}d��f�4����J�f2�,����Yq����%��*^��̷ߒ�x^DO
�8�����*��1��a��ЧQ�dNېiG��S}�\a�J��j��UB6_	/�Z��x�	�K��,#���l�-�[98C�DrŪ�\�p:��Z��q}��(�n\�G}2Q�v�,�4 \�Y�_�:����4�������^�?=���Y��i�>������@���f�<\$��,�t>����
vP���QxpF����j7�I��i�ҥY4���N�9�-������ʭ:�����Rq�=�2�ިĮ�QxJTs�2�~x��j���!)������C�����{\�z�^8	~�UtޒO6�[��P��G��aW`�ɴ7���MW�C�zH��Z�E�5�
�|�b�i���-^N��7�� z���Z�r.7i���ҹ�q0�91n�x�\(�N���yp6������_L��p����)�y~��H&Nxr9��ܺ�m�|�ǣֈd���٤_���U����R>ޯC�~��7�B�Y�q���|�"
�z}Kv�[A�?�<�a�������<�����Nɴ
O����Uh?�^��1���WcG�R�N����bJ�����|	KN���\�&�4��#�$���9:���21+&��y0��D������j~�Ι�N@,zn��Z��X�����P�7�X�� �<#����ag���e���Sn�/��7
���Ϯ�_8�"ЧQ��|t%ڿ������`:in��+D����%���&$��Ɉ7��EO���ӆq�q��ql9�^9�Έ�P����KO���dx�lH��H2�59A�����&ɮ�v@�\�z�׾��cv&7b���P����A���U��8�al��6���
 .��'o ���y2#8Yg�&���D��ӤaJ&��~!�6�n��P�Ӗ$a�g{���]��/���C}�h��W|��������r)�A�#��,A2�>B��{*��+����'��0�m���?֘�A#����:�0�Ґ�6M�Vl�M�A�n�J~
18#vHn�Hq�>!D�c�g3��f1N3z�5�Pv�-��z�j���R�]9M�[��Wi��ͺ:A�6�h���#�el�`m«��aP�J/ ���������0�N��)޶:�k�)�6:�k�)^�N�u�רS<W�2Ѩ^�F��5��Q�xn�Zh�o�K�AX>0a0��&��e��ߒub��~ߏV��Vk��j~�t@	��S_��i�RӔ��L���h�C�61�C���/�P��O�!��]�ݖ�ޡ)!@z�DP]{��m���q"�X����W8�����ƅ5N�oxi��y}��@,c��j#J�r��'��:,���d	O�&M�b��(�,��N���q���4'!��MU{�ΰm+p�L(���%nE�H/p���2�2m#Z���R(��� �H�h���ʹ�a{~�v��6�C/��,�u���r�?�Y���5���Sǁ���<ux���u���Sw{��<u]x:t��Ё���y:t��Ѕ�#��x:ڞ�#��\xz���{��o��{�޻�����<}؞�<}p��Ox��=Ox����A8p؟�����x�흖�i �dn�t�X��ݘ�8�O�<u����Sǅ��O]�����u���ӡO�<n�ӡO�.<9�t�����<9�t���{��;��~{��;��ޅ�<}p����<}p��Ox������y�����F�
/,m%�YSA�;�
�W~�C�X�����r��(�����2���O���`����>������bP���To�A�Z��4�;��|/��I?�DF����2�\�/��Y��S+'�`pA��k��7�%��'�qڏ2��toF�C�N��r��B��J ����|�>�/h��(Z�5�F,�z�s����L�����ѫ�+����z��+��#
J4>_���7Ǣ��M�ӄ��h�i����2K�g�d9���+�U�N��:E;�]���JH�3��A;K�|�I`��^�N^ɿ_�����g�����ձҐ�7�K�S���L����������P�7��?+��Y����o����������}�8T���#�����B�}�5�zC��c1-�(�g��S��\k�Roh]"~U�߯�߿�������5����S����������I �B������]��M1�!�{Y.^��"z�X/Q3�3Y�%�^���T�}��b�ŧ��4�H�7=ı�bNV�~��y�i3��~�)E9�kG�+]�od���9�(J��t����*"^fx��,� �!�g��5s/�
�B��U=�/]M��XGY�>��h~�!��П�d:����h�O/�Ct2���!
&<Rl�B��D�.;�Ʃ��c* J���6�;��vk�]�koЀ^�W,�%���O�N��`XDE��h��h'>S��h��cV���N{��3#+>���(&���#~>]�g����8ߋ��Q}.n������=Ҋ�7��@������A`t�g�Q<u���i�F���	�M��h����";���Iۮ�\tzbcU�τ����}`[O�˝t�F��zdٿ!����~D4#�<��]���7&s+�Hd�?c[�.-t�����O�)|�S�llAwi�k���g1{A���b�Eץ+���ȁƑJB�qd��KA�i�P�e���D�.0g�;Lзe�X{Qz�st��.1�pJ�7Q� ����R�TeW��*���g
�~ȗ=Q��'
JG��c�b{*��EKK��+�b��2"�&�\�v�$1	��]b<��oS��=.�(�Y�2�N�[#Q�[8�� ���0�?��D#��o�E�5X���Sn�B�:I����������2W��T*`�ջ�����gϐr��z*�Ft��S��ڈ����H@�5�</��B{;�l�����e��;���w�]�*,���1��#65e���E���KŬ֍ȕ� '��4��]}�4q1MQ�C
�b�r��[-�'9v��-�"ǒϓ��B�8����U�h�*Ok-d�!a5!SyB�U�TI�Ȱ�((�|�X��\��ۑ���s(J��'5���[$�f���k�Z@l���~��s��E��~�Jn��D��ݮ�gɼ����D�e�6��$������Ɂ��c${�$G�� ��:@&7!���M��Y��^jL=㱥��o;5Lg����:=X� 'p# ���֑�f\Y���7�(r�,T��8ì�r�!�*m�8	V^t�2n�.rr16BV3� >����v���5U�&��(�w�!�v���^��6B�3L;�EK�hJ����^���(M�H��	W�%M��Bȭ�v'�5��f.��/x���f�1��IMQ��+d5�(�aׅ�jv�
c}@����%BO��w�MN��ik9sԾ6���8�͚ay-�9����#J�.��n5�9&}�A�Ä��&^���;X/��kR��zAz�����߹����thH����L�R2��8��{��3$��­OƏ����2@���Kf��fmrZ��Y��s}�r3XMM�F#h}s��z��-sC�dOM��1+)��J�`�p�����KJP� �׺k�Z�!�'�EW$����SDr8��0W���V�^��J�'�O���`��{��9�&�(������2�U@���"��Z� p�PkS	A��6�Mk���L �R��j��ք��5d��hcH{�h�;��S��ab��V���O�&nˉB/�����]d�U'��8�A�����\w�6��H�{R��LoY�l3%��"Mi'L�����Ȫ��̇�Z�28}-n�B��5� 5Uf����ך�X�Q���T�������o
\h?���Xӳ�f��<Zu�����)9Zu7AK1�!���Nh��E��`W�eU ���ί��Ӱ�5QxR� +�Ug�y���8�����h�z�0|�T�U>�Y>��\�Y�����B�YrYd�ڸ�4�.��3�
�F$�8�d����c����
�O�⌆�w%��SU�V�b�E9�	���>����≬t>�j�]c���2�Vx��oVfO�
��M�cS.LRzR6�L�2��T�F�Wv�d��p��
3�4�\C�i5nF��t��*!_� ���u�3�������^��rFaS^̡���"̇��K:RI� �,ja�e�-�;nG�V��}�>�W���9S��h��M��c��szn_c���,���n�de���di��F���a�r��9�FIg�v�q�b�D���+S���[���h.*fq�x��l���V�-�,���8��j��C����&�)�VQ���yQo��I{��W=�c��-"��8yn�������c9��R�T���DC���{.XEP(�,C%�����yFN�3�;w��	�m���H�7#r'lW�r��ѺX����
%20LZ��U�A��4I����y<��"�,U��?������$�-sd"y-��ܪ*tN�47?��g
�r�6�U9�H���ʆ}���5ʦJ�kӯBo�b*��#GEP+q���0�$R�[5��e�ￒϻ��A�b^����v3P*��6�'-b��|.un�(%#n�}@ԑ+D��y1z�=��J�,�X����`���3�S��rΔ�r�7���"so�ro O6h���yb����Jt@��j�bX�t��si`K�#J��D��v�m6�W/YZv

q��F�"?A��h�T�o4�j��LW�!�h׹+<���7�^t°ϐ�禍���)C'N%��\gՁ��y�S)x�!n#�vvj�:��JN]6iSVn���h��E2$N'�|Ԝ���Q̳C�\�9����HAX�%s�i��Ί��f���K~��zx���X�ۈz�Y�X�c^�tq�bw`pH�-�.(Rz�g���n�.��$˴�&P���e�x])zw��>�%\��5`8��4�^-�=-�o�Ls�LnD�ϧr��7aT\�Ƕ�)�מ'm�Q�1��l����,r���&�ܳ�\�
�v��SZ��c���;����%pDQdT��t��U�'��~]c&Y�_��~��(+T^�@���G*"�J�G�S�S#}𫊱�g��;���7��r�h����Wa�����P|��O'�����>Y�h�(�)[������RC�$����@OJ�}QzO�9�����4��є�V��ՆXBN�eE
s�@D�Q${�5��+�3��M>#��Z�E8ڢ]j�f��d�V�ݡ�C��$�PhWB��l�*H?��@��.�PP�Tw�7Jh���k�<����$�	h�ՄdWbt?fw���Ic�c�<�]�$×np��Ix}����պ���u�(PZ�Zm|c������`#��򭸨U��PJ�� JmyD).�(�����`H��f4x��x^�(~��������~�#�Z2R�s��>R� ��k�O�nP�?/jWW��:O����50�	�]�����:$W��v��ժ��V�Z��jW�]��v�����ծڗs�/��a�j4ۺ�6���;0�ևĠ�C�1�g�1�'����������O������P��f������՜t��<����b [��g�kc�[�zA��le��VX�l��VX�l�nVl:�*�S�?j:I��a2��ؔͮ
��UA�*�Ʈ
��UA+�*heW��`+�*heW[�UdW����L�z�(��2i4O�<շ�ڥ|��kx��?�w�mp�#���y��P�֮��yN�x������-��ϺK���w	����d��Y�d�������GY��,?���g��6�視�;��S���6>�+?6li�z��c3��)�Ӥˤc�te�lm:�3���0�ߋi�:k`�o�b8���D�J�u�.���`�p�ns�~#8X-GtF[���1 ��ep�X	� lN�Y4g����?㤦�y���ڜ��E{4>v��.y�:���{���qy"��-ّs�q��(���0� �� ZE�����x̙��w8�Tkp��ܱ	]�V�ҎHف������XUZ�Uu��F�@���ߥZE�	��9��S�aP�r�b��s��D1L�r�A���b: ����w~)UEib�©6,
�Wr�+�d�����D+��D��iUw` ���� &Z��/����\.��آ\vǨ��i$abrq#T�4)�=X/��J�s,,�Y��F3L�qUY�}��?\�����Zc�0���B ����[r�:1�W��ZZ
,�߀�?��Q/���u`�I�`�QO�0�	T�� �rt�_/� R���@�Z6�Aښ��N2s�r�yy�<����j��Z��or����
#6����f~��A�Ck��"P���j?�2&$��7�ЗJ=5=ϭ_�R�O��f���m>��M�Zj�y�ki���Z�)�� /�[��'������͔�ǳۆy�jF����h��	%l�xy�������LnNl���%�T��|x2',�Ic�<R��+o�QhoΉ �-iS@\�K�d��#	V �l�j2�Bl�`2��7o�~�/Ehճڸ*�Sڌf[��f�*���JV�q#Ss��Tq;Eu���U$�9�H	nvYT�Ln!�<Լ�b��$�J����[+`S����Z��L��%PO�7i�y�z��󛺦%�����~� +��ӝ�"���������=��{���|&���#P��>�p�-.��,a^Ή������c|�D�q�Ϛ��GKʵe~
����:��2��rFJ.��o���jEj�.J���g������R�^��{ޱ�$Z	�`����%�\�%3�锧��7�.+�FI�g)9�W�[H�'����Xx�A'z�)�"(��(��^�ڪ����e�r ��`�o �	Ys��]�@��Z`������ݶU8��P%��ߴ��D�	Ťv�ܻ���Zsدc4����&p ^��o �_�׬w3p���x�	��m������ `S>�u�Ŕ��R7e�л:��O
�<f?)n��y����rU����p�9 ��7�t�l3�����,�#c�rNY8�X/꺝6���t���j���&�p���`8�ގ �$W��Ś�	>Y�\\FZ���e��kOD�aM��!��@�W��h�e9xc��K\���"��@��"�N}��R�`�|��	�ʛ�x�J4�۪��%��9� SN��A0�k��G��ùb� �
�kAsU��T]F���p�oE]X�"�|w��������K��gvw�>>�]_���0u :� G���t�A��C2� tg	^Ԛ�D����kZ0���5��8t~��Ak�_�GUGВ��E�R����>UW�Kf����bg�"�nA���{��<Q`�iM�A�h�.��o`�����Ұ��[tn�F8�ZS�R�em���_yo�������2x��n9�����Ɂ-< ����轩<FP��1n�M+�&�#��ⱉC��h��TN�F?g�gE1Q�><9�_�=jJ􃢙,0��Bx%4o�z�9�	�Hz�|���>���'�a�Y��-y��e)���g\;������/Vh��Z4�\�/� ��6�Um*����Qz��^ɮ��"/�ZL�s�}� �[q�m�6��|���h�+/�h��H�y�=�cbvSPz�rӝ��4��L
D�m�U�pĲiKV6V5eF�/Mh�dBg�m���kHȵ3�n���Hov��h,��v�iE����\뺼#0����٨��Ĕ�	�8�	F.a����_��)�%ڱS+0�R�˥ЗK�/�R_�tK9Í�d��NӢ�2:a�=%��R�+aV�ADpJ��Y���!��{-��UL'�Ѡ��*�L�@���}����h���Z�����!���y�M��x�ʳCy��y
T�c�O]�y�W�r�=��\z���	L+�`S��i��a��f�п}T�=0��2��ĳF�!��0���`{�!p0�?p���ݜޯ�n臶2Q.u�\
E�T�r)�n��x�'R�s�RffV���M0��e��m����&y��m�x����n�/�~���m��Ӣ�"X�%~��1�����P��%~��L|��O|��O|��O|o[|�nP|��P|��R��W�W�F�Z����Ң�uƶF)eF��\m�Ė2�M&޳�,��u�`�T�Т�����A_�������?i�z��.��E5��*��ǋ���Y �Gh.T�Wcw|�u�3��{�O�4���`�L� Y?��b���k$}?Z�p��j���'�/W�
�7����NC��0xRiNn #��oy�9
��@�%���)��1%~��/�d��"�Z��j��њ[9��pW6Q���+�"2��=m�8�ŉ8�V��zA�9���m2ށ�ԍ�Hg�䁮�����U�+�F.�tX���-'kӵ�y	��'�+0@��_i4�P��k��R^��/�B�
C��ӈ�z���8\y~�9�#�\yO.��f��o�]��i0�#�l	�1s{��2�By�܌�qǖK:��Z�Ǽ��c\���j�C�KC*\*��lJ�k��+�.Lwu���,�M�V��*@k�Z���w)
�o|���g���C�h+�dz��3�Ǻi���@̮C��� t���8������-o�N 巻�ñc S��Q�@Ki�N�&��ϡ;bC����&���o�@@aD��^v*U4�]X�=M!b���!hԌ��Wz+�*���d��^pc]��B S�!���J0 m)�c��8B[J�����;�x�������\r�^p�^r~6�<�_�3�<����=شA�[Ol�9��o�yk~����`y��/Sw��M{0c7��#����r��]�U]��� ��S��L@����+�q�hg�g�L�?�+w�J�D�i;Ro��O��O����I�`�R���L�rj����<���	��K����f;�S�쭐�_�V��#����]IUͽ ��^�_�[z�o����4��;��gt��WY���q����Ug���U�U)Z�dj���!~�Ë$�Y�S�}v&_����hL�����eB�牦|�[�	S�{�R���Su�(&r0
;�9�:^��ӭ���So��H� M�"��iF{MM&+z�_r5�Y�ق�''w�^bRX&y�!J���~!sFh�R����4�#^d�f��_c7Z����7տ�}���7���,7�Rf�a����$:�'ѐ^\��$�7򌓨�@t:���Du�9L"1K�_�Qy~��þ�=-gwi������!]��ݧ����}8@:t(a#�=����>w�YB�MC�Dd��IB�.�b�$)�+��L�H��ǻ��K�]_1�eG�V��S\��Ff��z<]Z����b��G+{vB�*����K�[�S��&�x�i��{i���,�K��k{\C����=)n2���K\ϊ:�yGŗ|��w{`R�	���@-���-�����5U��F6�ڻ_%��R�ǝ���(��b�
%�M_^��N	*b��/VJPx�T�b�H�kA
4�Dj_�D�h#>:��Ī�jVML��iv�f�����XlxV37EB    c6d8    2154x��]�s�8��5_������#s㝭�M9�e�,{2�WS,Y�e]dQCIy�_x�t���T�]��B?�x4�h�����6��~�[r^܏�����FR���Z2�?$���,'�?�$wO����m�<Y'���|�>A�q����ԵX%�f;+��|1�o�M�%DkN+i�X^��ն���z��Z�
������?��+������j��P
$-��E��>�]��DS�j�E�1��NL�OZ�m9�}�<�>�m�j����N/�LK�n�z�U���Ã�m��Ӵ\o�*|���*�,�Y�~��+�ۺz(C���Ŷ��p-����KqU����"�-+���+duE8*��^�,1V��a�e�#.�����a�V��g���j���?w���O@��8��-�1��h��)q�T\5#��U=+ꃢ���d������V��4���@�,��]}@�GK#�&�G!��M��h`�b�/��ź�ݭ¾�5-%;KΌ�lV����zvԳSz~��{��u�׏��@_!�듴"�{�( ˕V��Rz��M޳g �:ӱuhi\�<hvyh�ZL�Ŧ��z\.�i�th��HZ�$>��%���g�J�ŘV�hU���3!/h��).��㤞 条�z��Gt�c:X%�F�[���͸ߔ��lu��;KK���u�ܕ���q���:��'��
Mo瓺��Z��SE��#���zR�a'r��r�ڰ�����������V�:QJ'�=ك�D��-f����[�V\ﶎ��Ks7,DU�i�al8-�\���?8I�����V�f���у\����D6̍������|��]��b#�R<���кT�\��B����b�<n#+ӱ�>��E|Eb��n���Z�C��ʏ�<XiZ����m1�-���XZtj3��/=� h�w]�A�h�*,��g�����CK�πH���O����ƣ�-b����h�b3a�k/m�Q!�E,��
���+D�>���o��I�qd����Hj���L��ȹ�a�V4��{���{h���wd��4�x�����沚�wkR:4������)`�}#ʠ�(ɚ������'d1�CК�L�5���ؼ�+7�bȎ��� dip�!��Z\�j�+wG�u�����8�����$�`�+�l
V�<��d��bV >J�����fcc=��筧�[#��{^S���f��{:z�UO�K&��=>�5r��+��5n��f[e�]���Â���<7�C�x������B�QK���o�]u_��i����=�I�&���8�'��S��ɳr9�4��H��Ä M:��a����r�R.�p]���qWO�l)tv�oӓ��1A���҇$3¸Y��Rp���ā	�9�~�@Fsyށ��Ï�b�O��eĝx���l�]`���='�8F���|�,�n�M���A�+��9��o���
Z�������������Z\�[ P�;��Ќ����p��Gm�XO���&Q $�p+JȔ�gcw>-f�0c-u,�!j���M�<�4��O�m�^��+Z
5�Sg3IK�Hɪ��j�=���(�W�R0p(A���wEXNNs��"��L_0���/�jP}�i�?+^A3���N1�ӝa�,�#�`vhP�:���\��u�,�ې�Ҵ��x���mi���b�����	�'���%�찮����G�R����f�%���_�˄��4�8��s�����F���Z@�-0|�.��s7�`��l����c��h�g��%�2/We����"��q��!@��2�%�&�]͎N�j�����O����ܾ�9��*�� ������ߋ��o� ���'��I�i�\�>�vYT��F�}1����wqy�N����zs������Zv��Z��,�U�v�p�� tu7����Q�B�-Kq��o�Û���
�e��J��jA[�ٞ��d�R��lp{;�tD�&�弬m���/.��f19퐶G������&>x����{���{��et�8_������D��)Q�V�;���2˚���ë���0�s��Tk�jw�_�c�
�!B�]���倻�Ǣ��8KqB)Y,���QYV�����a?"N��� ��C�d��`5C�BKu}Z]��P
�+ �%v=D��|,,���v� ~���"A_�� �K�	86�8�&�6�&��T0�%@�)DȈkέ,�R��S(t
���D ��f�@��%����(���8vsM�c��L���e� .�#�|�-
#�Q�(��3NI4�<�&����x�E~`
(�`Am
��<p��f��K劻�(·Q��f[#f1R6�(��I����V!
|���Ӿu�z]US`
ˁ#d�

Q�,;��!T�L
[�AK�裠%�$������"�s^��Kڴ��_#�k�]��^�����~���1ty���y��h�|�P(D������`
(���)���TPax�"��d��JD>���#�wb"��w'��F�����J��L�z
�����	C��HR3��3�0��	�"9H$��F�"M��0�P�@H��Q$�U���(�r#�?�:J���0D���/�6�(��>��%ԈF)D��!:���X4�#�c>�;���<�R�B �P ��z��\�?8w%q� 9^fe_����k�"���l�^�im���(�R�D��h����r0��8� >�����u���A�vW<ojᴔ��6(3��sK�w6�}ސ^^_*�= �ş��-�e���j��B��$'"Ԝ�BC��_t�_tB_t _t�^��^t@^t^t�]t�]tA]`����A
����\��w��_�gl��w�}�~;Y͸��c�(!�+���� =���az:To�O?Ν�~��7�1����ʋ3<n��ϊ뛳0�)�m��{�����[�͔�~"�P�c�-b�6*�p���u���_hW/h���3�ƈa������\�����a+ߤr��n�Мr��BG�N�����0$JC�j�| ���s����:�\��Y���Y=��y1_W�b5�;�0(mԻ�*�񧞳 ��$���+��dYhJ����=g8��	�-�Es!f��A:
��T�$�ŬL�r��4��c�(4����٢����Yq9B��c����÷Y�]�Ov>8;LBܒ(j���.��5v�Ӗ�u�=9mڛŋ�����V[��&ڷ2�e���7��,7�F�o^�ý�|�7��$�4����$�10�9��^L�lW&Q�S�)y0~7����h��VJ��ZV�����hS��p{���V� "�_@D4J���,�z�wT��t�Iz�gDP�M'q����Mi}�w4��ٴ�����F��܊C���������R��>=��qZN����cC���������苍�$�D}@"�0�W̦v�!��X̪�f��al���x��{�D��0����T���n̻�U����c�ڂS����X=��C�Vr5��^m���L�g@@]GR�Z�����,v�(A��D�um~��٦6)؜�L�F���H
�@�ſ����`f�� �07o\DN�m܅I��0�N5]N'.$��BN��������ֳ���y�|�ܵ���v�]�Y��9w��f�z�;$�%NY�܄���U5f�*�v�D�/Uk�����/������v4���RK�����s�j���u��`%u��\��ID�1ysh��}�C��p��ؙ� 01shbb�g��900�ד{d��?�s�r$��ɘC����b��8?0s�HD�e���T3��ɂ�!k�Hm}K��E�a ��׋�cF����G�;�i�!��YB#�����Ծx��[dd�m�u��`&�1����X��)�'9�>��?��W������z#��#/ݔ�O��Ī��m7ߠ.�aE���[Ρ�@�;'N��{�	�@��V0�99W�\���`g� ���R��n2R߽:x��Sloqm�՜Վ�}Q!��������a_�x1?��}Oѕ�A	�u\��*�d߫:�*�cU�uVnMS�oz�ī�5Μ�f�F�E�HgCU� �Z������ǧr�Q�r�.�o5o�J6�لx.�y�LT1��U]�.��Ʉ���v���J���W����l�bq���x-FCf�1�x]Wb�w<���%^��r�X)�LJy��(,>{��S�s�P�8��&���Ψ'~��'�$��Y���'�R�į�0����,nw��p�����p��Ʃ�6�͉����FSm��o,1}b���f�ћqp�[��'������l�:^,� �Gn�_~�wzxgs+]>o���1�z�הd�3w6/��(�+��7�����\ͷO�ஆ���{,��@�^̟��S�Q֋��%�����2����0Vݧ�xߑl�,��#x��B�x��a����5��}<?���s+�.�=(ƟuS��|�D�v35 Z�E�@�[r����6����@�Px�1<<�_�#V��h4}`?�5��21G�}`�43��.������W犌/u���b�^�_�A�{2a��\ą��S�T0�%����d	� �mIq�$9�U�O �i��R��A�$�/cI����2s5�`�	%���h~y�A��HS�=U�㬎��Z'�L���^c�	

�� ɑqs?$X
���n���܉R#�4�I��Հ��`<T�I|!MB���o�R�L&�EYТ�nQF�(�[��-��et��0���瓘���^eStpe��.��YI`#HW/翺�o�������>	�ͤ��e=1@�e�ݒ��dD{�����u���o�����a;��)\{�%�?L4�!$��� z�^��hDn�Õ�?��S��F�z��K�t�3`�#��M��������S���͍Ӻ:[N�U��@0�?v�ɀ#�?�L��q"�k,�ު1����U-N�g�|�f��Q�G�+/o:y|8��"��Ǿ� ÄJx�sK�0m,-����b����Ҙ��jIi��d�Yl��ź��c�	�t�J�I�w𺉺b�\��x#<��r����3�Gir�sUv�{p��c�}).�����+�O[�z'5A�A&[f�kI�}�����'f.����4݇<i}-��I
�Xk�rN�	�0��PZ|��˼+�]�튄f�v�k����{�y<#N�B{Q�{rU%�|��=ǫm�)s�D^<Q����Al��l'��Y�ûo�ͷ�>����}
Fg���r[ΐ+T���n��V�n/��_��[v���r�Z��?M�z�P��f�P��^
*[��K��7v^=?��-V�L�� �*�*�=������VΌW���ߊ����q���Aq��r�c����G��k$�C�6������t��b�2�=��પ�ؓ��kz�/�i�1�-�窪�'��gV���j�S��vd�l�q*��j�UK�p	��z\��W�rH�
X߹7�7���WW�j�����D^w���X��ຊ�_�=��;X��s��s: �\ح*������[B_O���$X���⵮X��	���y_T5��+X����U`u�V�/����������<o��T`�}��+<�
�����W�+:�*:�*:�*:�*:�*:�*:�*:�+�o
��A���vg��V��.��a�f�������C���(?&�O���~�m�ȤB�@��4�&Ѥc�tB�^#$�0����"Q�c�pB^��
�Lզ&�~��<G-x�[��y���t��H���=̟�H��T��,�n���o�b�g��Լ�����۱�c;n�vҎ�u�����y�\��ݦ��J&��Y�Orn�¾�g��o����#���r?�u9�VW�&u7=�>��Ȇ�@���A�'� ����u�-�{v��{����W=�^��S��@�������;�|�q�#�w�;�|�q��w�{��^C>�(�'��d�i�����������������������lb�+�b0���z�����Y����v<���M�Cb�w�*:�ъ)EG��cZ���StB+:��`�^ӊN(E�1E?ъ^E�u�W=�N=�b�j���j���j���j���j���=�(��ӫnC��n*C�~��!�a7�!�Q��!�q7�!�I��!� VȍB�R˒S���X�	�:`e&8��Lp��� ����N�!�f�@�Z.���i�����2��~����0zD�Z/��9
(j���-���2g��$y���w��"��J�5�q��BtQ�����;�~�-OA�4߰��nL�إ�$�P��|�\.V�M��N@�E��ڥ@��z-.�C�?��賷y���Ad�O���z裧��9�Mn�h�Q�a�O_�I��Β7l|�P#ޗ�c�˘)�9i~
��a�sͷ�5%A�(
��ǆ�೓q��������	�EJ�>uP��g���}�ʑM��X�_y��=�>��do���/I�t)o�������s����3����j}�b,���t?�ӷa���v���oqi�_��f�3㝕�V�����k��䚩/���ӪC�]u��l�P~r�Z~�mz/��aƈ�`O�U��:mt�<�C�E�]��N[G���N左ޥ~���d���Q�
9W�E��M�h���U�Tv����$7��^>��$����KU��y��^������2��T��Һ�Aʣ�,)��@M�6Ƹ1�때���K��W1�S�^aJv���s��Y~7��t
�H'�V�~7f�W����E�K�p�1"�_��m���Fnp8w7�H���+_p�>�N����p�ju|��Z4�JC�$>@���}��@ڑH�/�p�䂏�E��<�I���)ed(I��"\�y�.�&��j�g�
������Hڞ�$�ا�*d��&A*�O���I�N�;�x��ɤ��'?�/}'�ԇ�KS�a�������[�'+w[�i��,E��.�3+����ax�����Z���ůi���I��	S���ן���j�x5BB�Ap;�����.�n���%4�G�!0q�Ĕ]��/AQڿ.�/섪���6�]hJǝ�k�6 %�RQ�1
�i
�Z�
�F�������@sc�찧��	(D	r���y�H�����_o��io����M�PBW@�,��S�x����/��t!�X�(��4Aˈ�h5�Hj0���±�5�52ש�ɥ�5�4���@�ں4t�a� ǣ���h��x������ڈ1�c�ɀ#k���0?F�֏�a~������'"�<R)4%Q�N��Dd/�D(9MK�y"��A�!���_r$���D��X淯w�Ɉ��GMH�%�+;.���I<�u�p�<ːon
u���'
��{U��囒R���
�e�X:94����ï�|�t�HC~G�a4T�wh����jjh62h͇���g�Z|��Rq`�W��|�l�rG��zT}�%�N3��[?q$����><����nJ�B�jM���$>�Ҹ��GY���~���2�Y�E�ϳ�����(J��i�r�D'R�L߯��K~�f9y�_�ps8��_i�Ǥ`��>�$�%w �th��jS�,��,IW��.Ǭ��1�\��g�}-�aF���>Ì�f}��3̾�g�Q>ì��0�|��|��3̺�3�g���g��>��K}��3�^�3�H�!B �k�82�IsNB���.�[���j��p� ���6��)��0���/pf���,�.݅̚Y��0��.̺�����-�	�ͷ�o�g��zCZz�Pa��HOBhpˍ����b�(��[��c~j9����J��H���2~]A7���֠Ad��=�hд���qDøA�=3�mP�৶t~���R[.��dY\��լy���X���_;@uhi��M�ʺ�Z|�}Q]�a,�����̡5��+ 
�K/�΀Q��������: �Q�I[V���.yI1��}�ESB�j��tbZ+T�����0Z��6���U�[9v#Ж��5�A�������&�k����ի�ȂT�����W�7�
��!�UQ����BQE5��&6zl�xI��T�t�JB �(�!�]R�eK��L[�Ð��|����6�i��Uࢰ
�����4�Ch^�j��B �<�MEd�</�i�z�<}^��V�H���&\�w�7�Ug�O�I=}b��Td��G7l��fc