XlxV37EB    3234     8fbx��Zmo�8�ί���J(�I��=خ�Q����=mu:E&qi�!A�a�����yi���CIc?c����5���T�M�g��m; ahژb�Ρ��;��Dڡ�tUmiڑ�#U�w�cR�8�hp?G{����j]�~@;������ Pߟ?�􎢯��x�dx�!�z��8 D�(	��>�%��ҏ�s�%��N�ɐ��g$�gN���*�>����9�سq`�����ϭ����.��J���<{Gzz����`����	����~aηǭ�)�d��'���̽hD>9!����P���@kjj��2)�NR�	Xs?H�K<s�)x��$�G�I[�Y���Q�L=����M���,׷�m��~�6��i;�7����j��yta`)& ~�/)~J<8�&����z� G6�u<b#�0'r��7W�/%h��;�"��S��f�g-� �cpVg����a�����b8�Ν9q�~~ f���.~ȉ��&���c5��I�ny�^���K6�YGI�=����R��o����Es\礭��%��C(��5���x��M�r���;t=����!�H|B�&�q5���F�����h�:X8h�~p96�7��|�������gי8x@�`0�V�A��aHm����ej���!v�L���1�3��(I�|v�����Ob.ۦ��X�V��O��Oc�i�+�^�(l�a%� '�$�*̖}s�~�Q���ٸ��n��U`x���0��	3�����F�ksp��4`�5�tNQ�؋�&�/���_���P��E ΐ��&���У'Z�� �X���jI,5Q?����\8#��� �H��ʸ�~C[���������hx��5�v-j�H���r�Vm>94kdsR	�T$��$��I�{���L�Y����P��J��	��X0\G���B�����Ŀ7Y~G�q��������8���Ia�������!��`^4qhln���wl�*��_�*<ը�ҕ7!� Cop��d��HZ��')�RTO��򢖴��UFq�����JF^T�dE���o&ԫ������M<�9c�R�IKFR�����x���,Y88�#W]��'J�ٌ��>_���9#I�tD\!M&��vI�O�5��O\Z�>�L<���O�S7W&2W�L��*b��jc�����u���=Ɵ[TKR��)�/I��+�O����0��\<!.#G�y�WX��H��*�l.W�`
����,�QA�}n�S� �k*E�$7;���d���t��y����A̾�ߐLh����;��@��=:��lf�(	�¡�s�N�[����0���?͊H_�]rK�MAA�2��Ck�$W�('O���@�v�x��<׊��oU���v�����Nf�˙Id�W`��jgKI�-g*�f*�1�Ǣ�k���Q��������Nfz\�zy6=�����c����3S�������+�D���;b>�9%�[Уx#!S�$���
�� ��ڻ��4��H����T��tVl>00�����	 G�z���4�'JcG�����z��\
�ʃOʀE�Q�W�5�nh|) [��}MJ�J(��t*C&�]nT�PI[Z �q	h�F�ݡRm�Pa�]]K�y��y,�t���\�)$�d�m'_v�]p-��i����<�"ړ,"�-��:l�7����M�ߒ���j��1��Z������c�������÷�J��dY�����01*�3�
�����A�4j��JI�S
K�r),!��RX�^�Vp-��i^$�e����La9��,�>���x�;��Vy�D9�D�91}�7ѣ󈜔��g�y�J��|�sE��E�h�1Q���Ca3v[�-:ן�i�Q�9"�-�{7	��(>\K���EѦ8�Ca�28��E�]) :�[Ȭ�/|l��N��kE��"��Grqy1�0����C�_�8e�;���f��ʖ=%	���a���<C>6NI�0�tEHV���D�f5^]�e@7q�'Y�h��.�&�� iJ,T�P���=�T+%tcO�	e��ܦ_��lxD�0*�����D���P󌰃�,�=j�X�!.5��Z�缄�-q��[�@/��++�c�n�%���[I�$u�Uҧ�N9_w�֑1�D�ww�z�[��#e���֯Q�d��$�-<�]�׶F�͚����봺��@�~�����הՐO}^R�(u%�bqCR��iB�")�����v���^�Y���Ŋ�%@��n6F<