XlxV37EB    10ff     49axڵW�o�8~��}�V@C�݇d�R�B/R����괊L��U�D��eu��HB t{*~(�g����f�6��{u�{>�\\՚��|�G.L�%�C�[�ɨ1�v�'�sz�n���s➝��'P�(E���K���M����W��	Th��DF�i�g���Ps��:ڱ* Љ��d㉆ƙxi�/�T.8P ��rNG-+�?.�=Ʃ S�|(q��|�R�Xd*0o���%U�d����4�t�eU���O�jʎ3����>���YN���'nF�.fz�<w0�%F�'&#�7u�n�i�v������J��'oɔ�1R[�M7�B�Y�H�ٜ��A�� \��mՏBQ�P���݀�z���#6?X}���j��ѿc3e�����TPɢ]��	�
�6+��O&��"�Ց�$�PMaJp�	
���t�ݒ3U��fRb9�@qQ<2A�J���2�xZ &,���ˬ71fNkf8:X;p&��k5�EB�i��f��.�q��c�4T�y�f��3��4$1^U�O�9�()v�Q�SL�|�-�l�PC̜�g�'p�$TFDт5GT)��Et�������&�04�(4��$i�����������{����w5Ά����n׫a�د�ң��c��������ToX$�!'�h8?'$)ps�e��ڭ�i�uC��)6M��w*ǵ��xgh5�'2M��'3}������e�
>�,��c�h6��fߊ��� \H?��ō�h��TyL����c�������o�݇��zJKs]���x�����n�g�3�ß��@�obߎx+�1�D`a��o����<������w�gt���V�չ���%^�g�M.^Ň%�f��0��@���{��IY|��sg&m��=�H��/�a���S��ό�[>�z�����z� m��[J:�@I�JrY��WJ���)j) �"hL����9���s-z
Q�nڄ�����:��i�H�<WT�Vd.��"�H�/���w�o\��6�(�K�O�A���)���MV�.9��)7I�3�0��T�,��Mrz	�aR�q~����8%I��.*6*��&����9cM���N��~�Fh6�o�^�S��h���79dP��^5�����\�����