XlxV37EB    2d39     8e3x��ZYo�H~ׯ(8,y,GR|d�8�cK	��FRf'�X4(�-5L5	�����ͫy[^kg���뫣��n���i�۰���p�de�}����5t���t��w��{=�������	�����Ɇ�F����M� @��=�O	\X���K~g&�O�q��	�M$�u����C���������+ڏt��Bl����0�c�j/^����=�t>ם��+^����6T�x�ox�#u�iT`Ǜkp�{K��'B��s�2�k��p᳛�y�+a�=�Wu��%�n�o��,��+� �;G���2b���o��d���b|���ה��p��t�ck
��.[p�t�P����S�e<TT���s �9[��~�����5�%�)� �.	��r�0��4�� �
��sz�8���l�r˧?�
%�X��J7�H�>y��~fn)��;�����ΰV3�u%��@	:k��̦���r�����ԟSl�p�.%��bg�Ov���g�K�̤U�BQ��cBn�u�`݃�{��m�Y�бD��Ԡh$�v=R��Y-��̡.�9��[�wۦ���T��Xu]Z�ո�^'��km��0@+�{L4K�ix3զ?�g�|z�������o^*L6st���p8h`~��]oNLk���ꦩ,r%���`%br�ǚ���)Y�N��U���|�E���<	�lG_�tx��7q<�X�������*`�P�FCT?�F�+r-�`n#. �l�/��|�u8���C�7�_kW?d1�;�+���p��u�����9�h��u�%^n��A�F�!9ľx��KTO�8�,��\��5�=\1� _	�2��<�s,�H�����g������B���Y���33��L��|)���	+�QG�\��ɱ#�^!�J�'�5|k�Լ,�����1�"�@(.����	�)�Ԟ��=7�G�}�v�՗�����2�=�G�[!"΍uM��0<�^p�!>/��}�
�k2���<`�;ߋ�(�(�i[ſЗ�8R.e�� ��|�
��u
�����;qz�K\C:�����y��h��z"�B&ӱv�U��R���0����kIpa�*	)\��\�Ҍs+AMZ�A�a\�'�;x w�����RP3@4��L�K#mt'v��U���x��xI.��9`�;ȼj��6%å���d�R�+�;dA!�*W�aiK�.h���L�ԟ�2u�tQ�L%?�+�����'5����e��-���f���#��|&#�!��M=�[5hZv��qbF�X�A!����Jt.��|RQn��F��\hG��x��,��	o�DI�@b[$���b�Q�� �A��4��M���|���u��B��q"E���R�؁�@��W�OAW=��Pq\8�,?���݉�حv/�<�")[�nL�#�+�4�ʔ�C
�]�8���L�0��k	0
�8�ԓ����Ijl�����������K��Id������E���M��+mQ�Ĳ)��wkbZx�Y�u6ll�>7�(,S,g�P�C�����264���$� ^�Y�G� �!2�T�� 4<���W˺W�z���Q ��j�:��CG���x\o�O��	�?���ǵ�U��zS_Vۋ����b�R����I��'E �֛�3X�*����]�f���/M>��g�6r�(?����[�/���ZN���X����Y��_�p��|v*� �]�dt���~��7E��`<�/[y�$�xAβ@�G	�.)��\�29���e2��Nlb�	�%��׾�_�@�)�J��Il8�E�Ҧ�:H�l�៩i��I}a>�݋"uj���yEw�Uԗ�@jj�N�6TR�%�Mz��Hϐ�����:-��f�,���B��YG��ݒrE���*u�+
�HQW���:�
%LK�R׺"��6j�����0�9���$Ny�45,r�,��9��%D� ^N�|P}���S�";#�q��z��`	�ԕLY	S�7eN�Y�H+:��5�F�r!��$��YN�3�.���l(q���2�Ҿ*��҅I��ޝea���R�J܎p�}ŷ7����-O�QF��:�䬜_'�rw�/�`���#��U�$�<�޶f��h���;�09��Fy�
�s�-�J䃂�r�[�I��44.]��60-ˎ��5wS+����/�VA�T���K���L�K�2�xh��q�[��!�ῲu��