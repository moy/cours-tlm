XlxV37EB    fa00    2b2fx��}s۶�����Ή�ʩHJNk7����3���No�}���m�V"U�r�3��?,~HH��s��t��],��X,���wp��9��������l����������a�}�0<�GQ��:����ћ�K����v��:@o�:���$����>fu:�We�G�з��a�:-�_����������~��Y�y����Kt2�#Q�2���)��D��Bo+?
��ǬBu��F�"��,�в,�e��I�e _�Y���}�e�}Q.�:+rT��- \�,��2�[��D�Eo���ͳi�W)�/��Fs@:s�|Aw)ZU�l�AoZ,3\3���(����h���_�rUV�$�Q]��1�r)U;=��=%�l&�L�4]`��OY��������ߏ���e���X��K`�BG<���5�%���y��@�e��f�w�ʧ�s	�
��Q�"�tZ��,�қ%xh?�i��Ɲb��Dc^��G��OX�fh?��j@E�����gL�r����PE�VJU��(�_�?�(j�[� ���s�U�	6D-�|:_�V�ո#�k_�����(��q��l�MMe�U�J+�'���<����DE��{���Lq}Um�������U$E=�^?�*ܲYVb#<ǖ�l�[G%��[��r�ݰ��XyQ���)��a��rٗF�9ez͘&9PI��6e\�-�ѓ�����e��{�)L�橋1����t�;������k/��|4�&�$#X��¢�
3��X�0]���w��ZLq�V����EZ�܄�m��pu�f�4O���>��9K�i�-A�(i����vp��9�?F�`��.W�;�q��`�u���Ǣ<��=xR����)�����7�qf�!��He�����~�z�x��#�TR!������0 *o�+��t���&��"��#!�����͋O���A���c��8�Xؕ��ю@���?�T��Y��7��}ޗ��p�CK
�_�����i�M�P)�i����}H���Ĳ�_�����|�F�ĳb��S����`oȧ#��*'�tU��:6Q1�Tś�;<WbU��-(�+
�2[�s�>���VG��9��U2q�7��U�]}���4��5��%��Z���T�/���Pf#�.W5"󁂗��fx��Yb�W2�]��0�*L�S[�9�3�Ò˩?�q�L�)��je�B�E�������͍޵�"5���F/�� 5�zsy{~���������߷/O޺�؛gw%^��7o���B����g�xȦq�^�U)�W}1�%{)]{cs�}�=*n�ۃf����-:ODP>&���8�����F_�)�+
��pyb'?a��({C������'�#�A�.�1��3?h<��u���G{�/Rc�bReXp�yM����5�r�Վ7HC� o>O�e��u�_eV�R,z� �e�)�5��R`�l��ҷ�e�'/�r�*w,�x��I|AU���)(XdSp�����(�7�3Du+	��{v��9�&��v���f܂�����_HWmw�=����p8D���l���7�;�g ��Vs�'��eO�π���{���ҷ��O�{~)�$�?\�n�A���������,�a�j��ύ�9�hd9n0�{Q��)��BBWO�� �r�'_�&|<��FQ�gb��wHk���Zn�,#��TNt+���$�����J�0�(��/~)�\I���)�Y�ww:ہ������m�����:+j�"B'�e �WhV|ʱ�2+��d-���(y�*�v�w�h,�f����6A;�&���H��*�������tY�Mt���,�Y
&�K����o������L�LFZW�����NX@� >����U3��I��v�GK�� �nN(^͐����Y|���.����lc.	��U�7����ˬli�ΦцiR�_bl+��kt�)��
s��?g��y����)#��lԼwI���Ck}��ƛck6���]�8�JƋ�V� )� ߃vyv{�F��¿I��B��,�*۸nɐ".��dZS���,�O�k��`��d�g|�.���f�!�����%���ORm�41��p�.�ٺ��m���+iKg�������Vj�I��DY,��3�DB������у���#�g�%:z�~��>�ѡW�55�6t���,���l��ۣ',>�<���k��K.�<�8���;�5Z���?�kC�Νޱ��=�������vu}�Ok�.6hޕ�E�li)�h �N �y��}��"ի���*hC������hE��P����.���2}h�,�8m�Q����{n ��?ۑZ%ڑF�H��H�V$�R����������p>�FQ<�����\`�*b��}8{^���%2B��2#g�Գ�c�`����v�\d2o�
'���ы��:ȁC�kG��c��}�j�d��wT�����'�����E0r@:#���~)P�B/�`��y"i5����6�=���}���ަW�HZM?�!�m��I�	�+$����I�)�B2t/�C�ku#C�����^ӡ�ѦW~HzM?� �����>r�^Hz���I��[#X��Ԣ������u���m�U�M�����
��@�{%ué�CZ�V9���^���|a-Z��^6�R�9�H]sN�9D�H]sN�9�=��朠s&x��5��3���H]sN�=~H]sN�=D~H]sN�=����朠{&x��5��3�e�	�g���~H]sN�ɜl0�(��[H<�Z�߉rG�0���$T`�/Q�����R��S���I݉��IWC��޵�pS��z�Yv��N|@r�n
Z�e�6���H�OA�:���s�Ly����o���I�׬6-�iMn$�4:���ZP�.M��Fa�M�ﳷ�ȓT%���M<ҶC��.�&0�o¶���O�&�'��J�����k� ��ʘ}S!p�:*�R� "�Ä㱛}b5<�4�Z)ـ[C
Vs�c_�i9�+u@�H�M��H��(��ɱE *��!Ef���u��b��a�!���
5,�D�X��%��bzR�����E��,��Ɔ､q�a���ʱ��:w]��0@ӕ��
2�� ��L-�m�≳�C;��vl)3��≻���]7)v�͔ �[�'z��G���H�+�)@7�2�| �t�U�4A�a�#+��2%�@�) j���uM)0AE�Tcp��j2�>���� �n��n���	v3v3v3z0u3u3u3�2Ö(�udĕs�\a�'٢��\�1&ka��N&W|ܬ#\��pm�µ����*Z��hm�Fks5Z��Q7W:J���YI��!a�Ĉ��hoH`k�E�}B7������8aے5p�g��ӂӬ��DD.]n�#� ���]���ϜxG��H;�n̼ޠ|�� P��=���U/�śY�c�!�<݉Q���@gx��	
J�}�Q��X@�]Pc'�����������PF���7����k}>�v��O���w���C�0���:Ǿ�${�]R.�$:nS��|Z9ԶZT�,\����EUew��GĹ��g�-M�X���tB�vB�u@��|��|��|��|D�Z���[��:���c��)����6�#, ?E+�bW���o��!����k�2�`�a(`lWO���Өw[�����h���-T:���ת��C4�s\B���jH��O7��r��"K��0�u����Nf����~邁�1�z�u� 5S�֣"�0],)�y���	�$Z,�g!��B`�Yl��:j��,�M�֩��|p����xi7�b�����wU$\ �X>0��� �`>� OK/�]U�ܤ~�p]��H�s�z�����k�m=�s������q!�w9�m��df�r�&0�{�N���~,S�)Վ`�YQ�kuq�����j�MD�Ǥ���!Ӟ~��* �&�<�\�B0�	�X�g�:�.����^f� ;OM�O�!ȀF$\-�kY���y��]f�m��Ɍ�20h2�m�4h23ބt>���0�Lr�dIcu�?i�A�y,V��o�n�/��=D�ūe
�v,�
�����@7)g^(H�Fv�G^�O����������� ��1�x*��CʂE��-����Fӏ���c�� �����Va��`���y�I��D�|f���T�d��j������b5�!]�N��(J2�T}ɧ�e���%���U�X<�ʹ�0��2�k)���%C�ꓺ|PSD�>������b��_��5%.:��{U9}{�@�F�	����$�[t�� �A�����c(�$�:}�>>#ߚ�>m���%H�Ȧ\d�* ��؆��.{��`�C�B�u�l���!�5�ɥ˻��q�Tᖮ�,!��H:$g���M�		(�3�r�|F��Q���hY>M)9��2[�L�0{,�'H�SgsRHr�Q��/�y:@Y���dh���,�%�2���?5y6k �{J>%,<��8�U��2��-C2��3��U���p��ÖdT>{����zI�&��H���E��%sE, i$Nztk��#�����72�@^���\)၏�G嬂�.2$Y��^"�?(d�=)$���$]2l�`+��AnF�N���Mѧ���^{ Yk�z7��qXX$=&��� ��DlFʒ���5>j���R���gm�ȱw��ۥ�]^^Ui�T��q`�љ�w#U'���k�˯��|}ZX��Kd�_*��vE6�|�u5؏��L)#�L~�*CN=[Wb<���gX
Bf\bl�P1M^y���&ە��O^z�+ȋO ʠ4~c4�`��M�-�Q��`KcT���1�E8i�p��G�'���K�;r���h�<�����T�̭(��KH�����蓻���{!�N�����"�Q��A���=�/eŇ�Gb��5�᲋"?��Gg�X-�����@����UJ��$��@����O`�?�����/vƈ����9�Yr>�^Pp�?��v.b��vNi��=��X�s����EY٠U���U���w��oA�A
�Ye;�ŕ��~�Hr
��79�9E�b�8ߘ�g��
i�h���.ɹ^9Z-�<^S��Ҹ��ɡ�K��pR�<��B�&�L��/e��oC����z�F��Y��p���cR���ى��d7z�:�`}]�jJ`�u�"Jߟ0��?��]=�/m��n��`����ɛ��ioKHO.���+�w!6�� f��d����L#���鉔�:н�P�-�CO�Zu3�e{-c��ϐ5��Nc���C�a�K@|�������(��i��y�ѱ[��
{�-7C?�	E��x�91�T��aǪ�<��ƞJC�!*�MGD�g�1g�7XC��S�s�)��9��Z��e�k��rZk�m��3�t�I	�e���4����x3�z� �"W��]�b������+>Nf���z�	����u#��)y_�t��c�,��L���y>����A�6M7���U"?�ҶP��-Nl�o;�2����,�K�p6ip6ip6i�l��٤��=�qo�u;,P� }K�*75��$�C�wz䌢��Er�V���m/���TI���kms��L�;qx���I�v宧���h��7x+���S�Z�f�J��ji������U�j�K����f���`���=J����c!C�K�� xmF^�RvYD�]����բE?���!�{3���L%����U(O�M�'�oO�AX��J@&]���'s����!���ý����2��I'�~]���u�eX*m���� ��^"!_'>,5D"��Qm%_��X�8�W@��T�9M�zp@�cF~6��ۑ��z��TC�L���%<���+�WR~��k]f��k���ʽY�7Q��%�s�3��5]��;�c�r��B�q�0Ǒ�lmly+@aH���R�D'~%�H����!��uB����7�ɩ�M�lb~������/7X�R�dB�Hn���M��nT�~q|�l�A��|"v��b��IyK��*�^3u�:�[�5�o���鬢�w 7Y5M		,e��n&� ?e����)�"�\� 7�������tτtǷ�ʫ!@�	U�kRm<%,[�˳l��4A�]�(����
�����?@&�o�MҀ��i�uӣY���SxB�@�4�����#�Cy���$��#�t�g�.�۲��Y�h��F�;�3\ǜ�j�G����\7q\��){�	��܆����]`�9�l#�ב6&r�K�n?�������O�+�⌘|����$�9�L.�v�ؚee~�v5�M�(��­iD�x��j"�zA߸��G��z�n��`=��m\���)Ml��x!�c�x"w�e�R~j[�D�H3N(�3�y!Fd1;�rؓe�؄].Us��rNh�h�z�{�	�ߕ�r�g�;�ɝ>�ܙN����)5L�Tl��`��]yjS�iͳzۡ��1�g!UeJ�X�<��{�����/}��: 97�¾J��E>ڐ�H#�"?ސ�a�1�¯>�B2�3�B2Ԟ3�B2��3�B2�6CV�|@"��O�~�a�a��H���+��H
��q_	-]��.r��*�S�`�!��P���UAmXA8j��諏��٣)z�h��=�����Qs4E���h�Ѥ�� zGv��5V�q���-������B�h�a5��xU��� ē�)_�7�<A�$V��uy�fC����{���I�3&�;�7`�&U����eoI[!S�`=1�����6lU�����~�3��Z�|��딧��%ƛH�:X_)�ߘ�"��f:&���3�Mf�a�*>�۫t!gJ���q�t�z��6�<ӝI%�o�z��N��=��4�_�=K�O·���n8=�����'FwS����b��.t;�����ϯ�?^�\�2D�Ca�.2��E
����G|�ؕ�C@lnX�u��Ո<�&��$�Ml�HQ�&*����ڧ>���~yX%�lPB��59�з��=����Q{�*V"���-��Q';���=��'7~��^ �g��%v��p$	k�&����O�
��Q�f/Ą�1�L���	]�D��gM::��/���a�ې�&Ҹ��%c�3DK|��Lw�
8�Yku���,/�~KK���mq�[�p�4��<���>�Po�e����W.kg�b"�u�{��5Ώ:��c���;��|�hځ�gV!ȅ�����R� ��~Yb\ȿY�R_1���H�|��јz��Bft��hfm��N���R.���O�X[�t��������O���k5v{�$��\�q^���4E���:X��B�x�絁?Bdcï��Cγl��^tF��5N9����ʲ�0dx4�(9� 0�(�[f����r/u�^nQ��BKU�H�G�ʴ[T?ʔ�̕�,�-"�o��|ܾ*5�!U�O4�g����'�ǳ룯����B0#%IX��U�6ġ�r#��Oԙ���^C߶g�lC�~W9yv��:�j]Ĕ	���B��MFz��ښ�yo�הn�q���.�ԟ��w��Ɨ+�����zc4��9��C�G���2/����5$��������;K뽵�?��� >|(��4�ӎ��@��5(�j���B��EY�Ӛ�� +��<y��w)*��Jg�� �>fZ޲���*n��d��¶��h��i��B���$��7y�]��b�d+pn��I@re��6��s�Í�
�(��-����X���)�&�%wJȑ-\�f��7�e��Q�Q{������żF̆��#���
��?��dw�Pю�W;�5�#ܮv����nE;"O�	�hh�D�"���vD�Վ�?\;��h�hM�1ZWKFkj�h�Z2�ג��Ğ-C=2�4*�{�8mT�m9kT�킊��F�P�<+4�x	���0��eʔ�B+l��Fm�#�������V��&�G^�l��+M����Tv��A��|�o��J96��2�v�C�^��X���U�n�JsJ��B�?=�G�y��I%.�����̐r�ج�H^�XՍ�7s���ۛMX�K���Sn�Tŗs;�|0���͕�L���`9L��t��\�@$��7J'l��x������Vj�(:�G��b������52���9{�3Z�$@#$��X��A����&I�x�ީ"��^�Hy�/�$h��9��$hz�}G0��n)��Mr��[	]�2r�y'@�Z�� ��2���]���R�h�]�r}�ծ^�с��gx򠶅?�I�q��J�;�(l.^�������OIPJ_����R���y{+�!84`!�����V6γ��C�c����QNz���#7f>�y��L��;��������������5]5�Ţ���"B�:Ex�T����S�O!K5���U��)ó�#�3M���}{F{	� l��۷�ᰖg��,턡R��������VO�Tq�ˈ�E��!U��8��3!owf¡-C��XZޑSI�[>(^d6��v�¤�?�J�=��TJ�%��Z��³�e�q��N�k��<�^7�k��Z뺗�5E��yۇ�[�-��t�����ʱ˅{{+Xw�v�ѹ�h��|���rgJҿ���x���ʌk����;a�Hl��/*vO�ӍIT4�ܳ���eI�-wJ�f�aKHN��rZ��pҋ=�5�_����\Ӭ��ަy���5���Fd}�ĖK���d��(�H���`��1b7dx�ybģ��-�����A�7��6J�i�6Q5u��-?���	�0�
CD÷��3��^�#�#��Bm�P��L�̃�`G1�쐧I��|�=&�%��z`-�?����#�6b�(v���ϯQ�r���<���|��79�u�x��.�~ߙkѻ-f��J���!���S�ul����5{׳s(at���҇�v��q�] p�o�>�i��bK�"_�b͈�Qnd�i��'X�a��^�f��F��
y޶bYg���W�f x��=V��P��j��cʼl �(S�Q�5x1V&�7LL=�!i��ɤ���9f��R��1MN^$Ƅ廿[�V䘄=�(��"��h���;��
�q����k:BMR��8B:�VG�tR2!Y��?��F�@���\>0*l����ZO5�@�$��:��j�x.����k;@� {Jm<vV���<�#�����"O���P����F��$��:�����D���<"9�����=���q�� }�<�Cc~��������J�+�_�*�����'���%qe�p=���[��6`u��]t��m��x�It3��%b=�'�c��_q����7�;��<���!�Y#;"�^'���7J:m���n�����u�dz��Gu�z�j������ጟ����B�lӅ&�:�_{���K�4Vs�� �}�����mR8sP�aGNC���_[�B���v�
��`�]�|���*>SŪt>�0�~:�M �� �Y5��7"S�@_��MDL���!Օ��ʡЕС+v}����P�l�5�E���QՆ�P	��)r̓pm�|�˹K8��L�N�ȃzhz���,�Ot�Vҹ	��oȞpP%�XF^k2���lL���_��g7�[&'Y[�%g�-��w�Cb����c��l7c���JI���H�DR|�&PX�'�ۀ�SrmY���e=6v�G�뱹c=j�G���葹�=67�q��lOx���� �]�gw�)$�4�(��8jC�}�}���p���+��+����|��펵ƫ�����o������S+�m��E�J�7J��)+0��~��92VY�(%yz�(Hj
�}���=�_��]�o�"�\�e絘�^�	��k��/Ǎ�&&�ぞ"���fGj����*4w3��;�8��|Zs`���`���9b;[�0p��ш\�|�z:��2Y�'L|��֎V��DH�J� E��N5��V�
�X�c��{V~c2�M��硖����S��~%['�$/Þ�&���"Kvӹ�:,��z�.����f�c��8jc����l��p���n�F��UV ��F<<�Q�LU���l���m�:]B�-	��d�<�Y8��*��b�@� �pu:�0�����
a��N+�+�0@�oh�!�2e���	{~y~�Kٗ����nU�������F���[ܺyr�WY����]Ȇ�������2'RF~F�a��g�e�<��C��50���j�a�|��>� ���q{�ŕe`�eQ�M�����#���X>�U��e p}2>�<�#�W�!m�Hk �.��P�آ>��3��r�zY���چV���v M�Zvc*�������1�]]��.J؈��D���%#�j\e�㎔\$X'��q]�L��f"�3�?����v�:����'���ޡ��{�>~�a���/��7^���l��=P��8��xM�M��y 2P�oU�(*L�͡�g�<��(�G�t���U>�x��>����������i���}�<��v.�U!�jФ��L򇔜�YB\+i:���*(�8r�4�:Y�(&3��CYn+��8&)v���~h��p~��q.K휻�)��Κ��!�0oR�G�;�(xa�0��X��	`tT����K	 ���<y���sK�g�U�.��X];������;�3��^:X�ͅY�;?�;�}K\��cs��0nm�گ~�zp,���kI�S���K����KŴ.lݝaݧl���s�n�{��z��["��F�,:,�9۫%�sB���\"��i�1Sm�Z;��KM$�t�C�St���� l]��XlxV37EB    189a     4fex��Xmo�8��_a��%�v+^��k�=�M���\7��}�X�$V��0�e��$�l���
������6xF�]���"�A���l��3���xMXe?�����I��>+��ar��D�b�6�L\i��<z���@t9�e�t��S�y��S�{NWl��re�Q�]�k��.��-���$���[H�9�@������0�%efpyw����`V|��b`i�S���k��6m$ŷU'����i�Vi5Z�r�`�,�:��j�V{�e��������G$#�1�L�%p� ����@<$�!#So����:�g�!{+��2ښ��-��ЋX�8J�_<�PN�y:(����5G�N��=i����
�^L�7)Af��,%�v������i�H2��y����U���$�9P�h����tl�ZE�#C�tʯ	���Hq ��o������~HI;��f��0��I�@�G��V����|�6Ux���$�Acv}̶��*)�}�`���F2oH���7<	���T�!@g��2�R�d8R��W?H�{����? �"
�|�>>J (���x��ɧ�I��
#�!�\�>U�� 6�´l�o&��(m����O�A�oI/ �G�ڈSqk#� ��ܓ0�����r�r���y/���/r@�‎� 3�c�)M��s������dK���H��L� �U�p��@T]h#
I�B~��GD+R�����{ �%��0����3��b�A��V����0ϲ���;"�He��R[l(�����R
V��a]M&�Ai\��]���(���)�+N;��*9����2i��4���}�ƮT1K\l�.��eHz_�k�Y�������ݐ[�@�i��� �^���KL_CR���g��ܫ�h�.c�͆9�ɨs9W%0t��_*�>�4�螲�r[����v��O�-2m��L���;�v�w9�b&�!�:�R�C����lKq��:�vֵ��r}NU��]-AMga
�K�4k�o�Y2�]�c��t)�M�]ʭ�U��8{��4������յ[j��Fi���2W��S(7�'W~���C_�),M�3`sEEL�w�ౚ�tͰ��p���;�\i�no��e~v4r�خ�0K�ݑ�5������u( ��s�F�+E�mAu�BuZP��P�T{/T��ꂪ���_DcR�U�S�����t����3�ZI�M@-g�*�z�֋�5���ID���=X�4��