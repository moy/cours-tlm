XlxV37EB    2eb6     b73x���n�8��_A�$�8��v��i
8��
�&��t�.�,юPY2(�V���9�H��ųh�f[<�;I��N컛[˹����u�k�G~��Y&�atq�y�;�;�~��ǻn�]����>�I��M���ڭ�o�!̗���9%4J�t��e�s�R/]3J^�#2-=o�2�W{,�S�-�h�!v䝑z�a��F�6�?�+��H��� ����)�$����$�#�L6��n�ť+�x,X�j�^�B��&$}��fn���Ju_C�I��<�����T�5���s�rs�E��W>�!b���k�	�;�?�����KRi�W��]�"9�`��Q2Pfr�4�P�[�����z��:ё�����ь ����Q��q�`�F~~�;�=�Y�B,��Ȓ�/hDY�5�
���VC[Cn�΃��$ݯh��ӧKÄr�R�t��E�Dt��W�
�%�xޚ1pG*�y:�/gA�B(n�`(ċ��*Xѐ�30��K�9t�@���B�䓣�^��-��YH��QP��� ����I�NW딬bhK^�s��&�((5�� F7�|1Z��C2�Ed���q���s�Qc�G���D�xߏ���t�*�0@�ԅ�tE��?ZwS{��|���o�s�x7���KE+f�e{b[�uނ�Β�w�xxN���37�s�/���Y�������:��,�?�.�+{2t^�bjfL_�8>`���]&L���*F5IK-r��],�IU)�/G0�o��
�/��������s��b�b�R��N<�gt��F�$)Î�?�r���Q�(#y5����ݒ$�>���I�}�\�0���}7���~E�D���ַ��0���& ?��b5��Pb(Gi#&/¦��|�
`A|�_ɈBh��_FRg�2�ke+�����ݚ0����t�p�E8��U�`�tl��l��I�ʊ�@UP�:���a�2W߄k���y�|Mri@urY�e� ����)����w�����s�w�S7¡H�b,f��ݯzź_��l`��-�Nye�nxB�p��N��z���ڒA�u �n��H�Q���Bv TYXh�D�G&/�I����u*�P�z&�WL޿��\���4Zh5�|,�P�� ���:j���>��=����8_�V����G���joS��ז`Y�1t*�P�߯n��u �fIZ�� ���W�U�@����M�(�5�}a&i��V}OKw��"
���̂4�!�C-J�t�5P���ĘB�E$R�P�A�P�Y$9_G<�������NL�H���+���b�n�y@Ԓ;<NV�.�Le�V�Y�G�si�
�R١��SG���r�	�S3�W�<{����~�<�f�-TVX�=�ѩ�5J�3�j"BIL�t��+�P�6�t��e�,�[b������*H�>�n�Ķ}��%�[�	��,���d9@�U�9(::SE_�sɓF�����Y�5Y_�mC�r���������~�/��R��9�s��� #5�6�����wL�P!��_��Tө��s:Y����)�N'C�v������)�I��^ ��=T�0ޖu�㧢��PA�
��-������&I��e��@�����h�h	ŉ�L������L+��uI
:��hI��-u���im�أ�賅N�����P0�?��J�=�	s~����\>9߭�=G�6��uVn꾠�աJ]�+���@QؚU6a>BX��B�ū�U��������_����*v�F`D5S�,o}�X�d)�X�.V!]�0"�Yr �..�$�S�[xW�6��Z�㓃�r�j�v(1�g��c�&9Q[�Nq���=:���h>��A�AN��t�g��X"�~G��-w?��|Z�:(�FjR1$�MR�Yg	xe����2Bq��N�e��	~��Yy���M���Ð��'��Y�N�1�j����Ά
��'����0�8����ԕ�]�[���K���O��Ҵ^�U���.e�B1���
�F�)�3��ǐ���Wa�a-X�lAj�	�7P�vJ�`^6e�j�	b�~��5�4\!�n�'�zF`s�i��3l��ג�Q�%!Ɗ����_ħ��B�eV(7]��M�,A�8[,)n#P�Q6}�h�a�$��"���L�ym�Cz�%��HU"r��S
Բxn�E�
�"UY�zJ-*DPU�F��Q���5��O)�c�u����'F�cf�<���e�P˪����@6��"���A4���\N���Y{���ߪ}��
�����P�J��:�x��hC�q�:h�H5#p~��%!-b��m�M���&j�uP���\�^��"7qFg��j�_Qn����}r���<����5�KS|1��y#z cT�l㬄��>&E֎��B?�~��n^e��g��E�t+�h��D�W���E���s�CSμfN�Z������'~0�S��C��H��Z`��^nF�$j{U��Q�����߄���mf�������ѿ$Y�=�����f���.����Y��#�Oq��q�-�L����3K~~i�(��#H�Ѕ<�]�V:�3~C���X^�,ݕ��0nF���c=�������^)�t3�h�M�oe�o�af�*\&������JI~Ò1�/�WNɿ����F\�d8�K�'����A�Z�����X��.�t�A�7P��OB�J���N�n��u��u�wK��M2�k���7/��K���5����{��S�'j���3��U�.7�U�'�QI�k�u�I *0;��KB�W1��	��|Y��uٯ��E�X��Q�3W��<��b�f�t@���+�?)�a�zU��8�����T���U�޴r��J_�I��q�c�㣸��_����f8�*