XlxV37EB    1b44     719xڵXmo�8�ί�+�T@!���`�ۥ�H�[Q����.2��VC�C�i���B��'�<c�x�;���u}yճ/,�v/+����>�`�m�t�BA�=fm,��Z�����Q�ud��4�''��)���!�z/3���%��\�j�N}���p�	�9���i��k�Ò� ��%g�G��c�K,�i�f@��@B܈��uj�W�������)m�kX�)���~"�V��$r�+�f"��3�NqgC�4�q5S�ջ0�V�
��� ?c���XEw.�z&'����|��KS� )٪7?֛'R���PĞ���ɔ�k!��a;qq[P��g��'^؆��ޡ��%(���r�F9��^M5�������^�_�2�5��SR6��?�>��)�j��}��͑���1�b9��->��2HL��`:�)��E�v��8g�9nGqN���	�#^��$.�f�36���/�	�f�,sj���&��Rr۞�:�8\�4#L�%`�P�����P��!���\�,�B���t6�.�C�H�|��2Y��έт?��=��3�p7�Qf����aH�i�e����no�[;|h� �N�	�
�ԻZ���e��yqw}���SE�c#N��^�ש A�S#���ح��q�x^fПO%�l�#��>sx0���^�ͦM4l��������db�	�4�d2%�
�ͅg�q2ŝ�B6�j��F��.�덌P�:�z��_�j�X��J%I~P��09��v�]����m��1��*,;
� 8=��|4;���;���s��}��[W*�)��� c=w��V�zB�e�Y��{��d-ޫl��+u�Ԫ�Y�=%Z�'2�F�����G��G��x贻��W����6�g��X٤��_+n�M�V*\j��F[�(W���z+R��in�����X��W�曡�cX�Pڝ�𴛽~����;S5wɱ�7���UiM��/LHp���#C�"w���$�N(OG�7�D̎im|������-'�i�f������ZF�Xb3+sV2(��B	�PI�����`#�n4�U�݌7�S��+��#�1����{RHMt�G]/1��Eۤ�EsxxW���,�����g��?�}F�.��/lb��^��@����{x:Oo��Z�y'��!���B��e@��'����qA_��d��-7�:8K4������H��h�W�S�ZU�#n�Qc��|�c�'M?jLݙm�[F����ԝ�ǚIӏSwf�5����+�r3��iژ�3mN��9y�|Tꀼ��5?�|ψWAi_�\ve&C5I�Gg0^:��EQ%�wI}L?US���$I��"u�}�i�<~=#�V)�:l�zdD=I¨謤rC��
pk����HT��d�T�\;��<�r�Q���K*���w�J<U�A�2��Z��C�ס���FP�J=ɰ��kv��Pb��Z�NY����O%ד��Qo�2H�V�|�V� �)�J�V���fN��*J-��6�g
'�'oUt}�|���|��R̚��f�˷�� 30c��� BVܘNY��8KY]Zh�Ƴ	�J�V�9`53�&�6�K���3��${	�d��72�!�_��rԶF�&�ov� k3��2���P�4_$� ��a	U��(h��dħ��� �D� �ʯ��(K
��A�@|�㜩�}�r'4�}��$fY�m9eUvt8��}��VS�����X�$*dH�q��}��,�TV�f��t)	�c�r�
��g(��s�`�v6�����ޞ����q