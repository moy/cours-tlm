XlxV37EB    2552     9d3x��Z{O�:����b���)Lۋ�j�0R��K��v����Z�Id'FW���9��8iZ��F#(�y�<~�8��ݑsyv>tO�1�5v��y����{˹�^��^��:��/�ޗ_�����w~#2�RR���cL~�C��K�<}��yI*�hC�+�Άg9��'�g�����	�=��aD1H"�db��=���>"�<`!]�~f�I���Ga�E�ݽN���	���q�o;�8`�$ɜ���-����4���9��$fb��"�u��/B��C��T	���ፑR	I��
*���>:��	O�GX7H�y$�p�Y$h�;�s�D⩯LS�9Mw���.�x77������&����3ߨ\���NH��S!�\�,#�⁜T2�I=�I�h3�J>��@�vΧ�D3�E䧁Ύ��Skc�����K���L�Aq$%��$����T����R�f�	��3�L&�ٔ��3�$T�X�N�O�Jf,d�JC�yA�t b�=mmf�S�HL�{:{�St�@��@�dn����#�}��E�FnC��E��)|�R�g�3��p�-0���%U!%A���OꞭ7�ʹ� ��73h./��j�_�ϗ��ϟ�
�@�O^"*�/���7���U��;�@�My�iy������	?aP5ІC(Z���~���Z>/�j��<�ϋR -��Q�-,Ƙ�,P��y���Ч�`�?��!R>��/Lv�iՃ��e�>�ڰΒhJ�4�S�$�,>^h�ْC����6����v�|6[��r �&๐< ��Д=
�]H�Ǥd�I3�o����Q9�qb`�P�Th����r������ӟ������*�
]��lM�iO&��6n��u`���V�Dz'�r�=M����}��q�f[]�SKGj�
�I�X�F���	bOL>�e(�cw��w��sXlF�'Cr솊⏫�Ҽ�x����ǃ���:��&?=0���1�{��0��v���%�O@�6��)�me����1���n��r�Qw�kU �����Mpc�7�	T�.�|��^3�U\�A�$�#��ߚ�?���I�\6�A�R�e�0�i�T��g�t�ʯ��H~��"t}�?�����Nu��9l,�lAɣ��+�����F&�������TP�A�� /T{-���ҜB�G��BV�R&q��%�hv��ݖ1��
(J�_��D��q��Zn��|�㿊��Zc�g7��*/���i� +4�W�T��˫�F��$M�U=��-��T��^�=�
���Cz��H�AÁ�ցH���_����\\#��ml(*��b���b"�thJ�T�u�{����u���ޏ{yagu]l�Fc����$��(�)LI�ИL�������c��f���D5 �JX%�Ip�����*�����J-��7ٔ��&��d�:킫4�#R��*]IS��"�/E�'�7��3��>I�N��L�zFC��HE���V�DWM#�)i�E��܌�[������<)+(L;{O�0�̨У^�,���'�A�u��v�ȷü*Lwp�������=^�c`�!&\	ԉ=��N�0sQ�[#��뀴�NX ���NKf��3j󹑿3 ��q;�<����.Q�8	g,qq�t��i+e��i�U���0��(�A��$��6W���N�Z�%�����2A��@�t�!鴬�Ⳃ����U�m{���mї��a������W��m�/�5�녵�e�z����n�];�W�p`/��P�x`-�Ȃ2��#���Se Ƕ�rs 	za���}賅v=}�e�|�`��1��>���Z�#8�@Śp��
d�tt�(�0��Y�mM�-���s�P}��aV�ӱr�Kz�8%5#@u!�5۝m3y�ڹ .�oY &z�w���i�xLҬ��X���׮�����,����Xw��[�
s�����S��Ye��YW��z\!L�Ҽb��\8?�� �1dEK5���U�A@3�ワH��5��b�Kp���l!�@�B��o�����v*Xkn��!mLѭj��h�Z{��ަ���vTR�Z��Y���<�\���l+�K���q�u�m����o�Z65&Gڕ��9�A-��Z驕y�c�)iE�
˿*E���v��	(S�y��
��) U�֚p\8��x�p�I@vUP����/���.>a�`�^$�]R���M��du�*ũh a��������d�Oy�!����3�\ R�&w U�0����i�j���E]���<
��.>�����ϫة��o��P��>�.d�t;|ݢ7����F`���}�&�̅�����f�V����[�|�ᗒ��]�������Q�】}��Ϙ��|*+qY��@>��\Da�J�5c�|�9��i�l:�jG��@b���XW[P�ϯ#�*{���	23���9���l�~YX}���&���