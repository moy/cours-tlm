XlxV37EB    6cf5    1284x��]mo�8��_AdW��f-%�.�@��]����K�p���ʒ!�y)���)J$E�Jjo��Ʀf���p�pHq߽.>���� ��|�y���#?��$\���NL}:I�����=��>��~������@���v�����n�H�qI~ކB��.#�yGh�x�ӯn4�{	�"��z����mŧ��t��S���	��|/xl�A0�#�'�OCL"��N�ؓ�����{>�=:����Q�AFEv��G�4�D�2��΍��ܛ̅��$!��d�)�#��)�8�Vd5�c���yj���>P��:�^��yv=�'��}�\E��K�{ڬ�{�R�������O���z��M'�dF���Y��'xqFO�\iVL0�Y������Eq"|vK
^�/�AD�1��A|��ѝ�i�>�؛�ͺ��	v3��N�V3p���u���8S��'�����ܡ1�$u���P �]r�h�M�X9�y+����Ȕ�y��iI�[>�rՓ8��M(Y�0��1�E��ť|�UAwX�o"�M�ŭ��J��W
�ĸ���g�(��#k��>)b�q��R�*@�u}��v$ou�� }��*fT�J�yX�{>HxG�U�\%dF����M�7��Ƞ��hd��̵ނ�G�a.�yy�9�^B$��1��E��1]'Ը^v{��ڵ�0@7�	ƅ����3�.ƃ����9��?���Ǎ��߻���z�^g��'S�g�ı�{��K��G�D�I&�ܛD��~�����n;.g+�ﱢO�h0:�k�&�M+�.#w�p�#�N��Nxw�isx���b�w�ifv���Й�tЕw�滐�T�z�N'Ic'�'G�7�EOV�uNO�'�h����Cqg��q3J}8 ��d���ާ��N����Y�yp<� ~��i��Q���t{W����Xn�Ч8=�,����տ�v��)W�u�'c�?���c���������a���;#I�H�k���pɡ�n�� �;����뫱srz:���f��+�ֻ;��眤��o�u�ۻ���Xd������$���!��ٓ��`��˾s��p����rN��Մ:�`�0j��%g}g5E}3�E�������W���z�R���� 5�t��ϒ']u��~NP_�ލ6[��s�E�0�-�+)�YU"]�lLQB0v�R�����UL([c�p��V��@ �w�a��FS�X�D`	�'�Z+��uL��`�Y�@��X��� ��uU/�]�y4R��թ8�!�<��$o�o����]6 �ޘ ������ꏰWp�R#�lL��s24®*^� =K����0�:��D��@x��N��J�3��F���1EnA��� ��:[�6'RZ��T$J6�n���_�B�uv*��p�|�'/�I:P2 �j�_��`QNuS�J�2�ȉԹ��43��+p��8��Uȱ�\F��T�_^�A�D$4α���R1�����������Y���S�tČ)y:.%�"�J��q�Q)Ӏ�bJir,SU[>�ѩ0;�����DRP*�bKyG�4!<3�(ʀ=����4��F3S*I� T&�`l��t42�h�D���t��'�]�D"y�a�pc=�]���R����VU��X�cl�9�m��ij!����h���4�6F,�:�����fK���x&Sb�Q��:m��5�k1��Ӄ�2T�"�����6B믘����F�СL
��D�4NBxs�M�򨽍�*Ss���-̉�{2rr�%��o0I��9&E[�R�O	2I�Q���ĢȻU��Y�(�#�.$3��3�(���\ǻ#=��ĝ�`G�0�Bw3(��y�0Nxw"b*�G��'ө�����l���'ƚX��,{ �3�Vw�wX7q/ؤ�t��b5������~?d�c�#�'��`!�a���D��ȁ�y�W6��� 2�u�d�TV
M�D�+��Vl�����}c��8�oR:�7[FA����IS��!72Ʀd0��id�`X�Q�ͨ7o�-���t"�s������<AR.G��y~��X��M�Gǹ�ևw2������6�V|���K^O���h��T���M�����H�Ne���E���	�ef�tU��1�Ϛ|��&�$n��v�P�򊙇�4�wAQ1�!�IaFf��l��\��֝N#l|t��O�`��X�KiA��)���u XWM��C �m�m��!�r%�L�ՔƄ��Q�b��9~�c��
!�<��۹1 Wݷٸ�����E�$��>��%zS�S?6(@�!��[
x.�r+Is�xG:���s�2�Tdv`X��FmH� �g�8óKx�9eK�JM]�M���g�3$�X[X�NlH�X�4��)# b�e�0d�Xy��ɐ;&�/�IY#�^�\g2d������K!������TV�m��%����0k&`f%�Z�Z�	��������9-�.�f�RU�KӒ��Z��9+Yì�����z��VsY���j+x�� rV����sԔv�(i�e���J���]�Y�f�j�5�s�5�Z��E�f3���fua��01k):`�JZu���Y�ZkkI=`VKZk��l�`�JZ5ji��fV�n��A`�aL�*v-jͬ�`��*��miCJ�e�v��~����N���*n��p��X��i��.�=��L@^�)q� ��-|��d��ݔ���Xѩ�.�	CR�>����*�{�r�Pn;PG��	|Ev���ٽ"�Wd���~(�K1R��̞*�:�֔xEv��D���n9s���p|�g7M��t��˶�q�-ee���E�h���:�����َ�/��M���W�l�j�Ӟ�Տ���*N;-)F7�	1B���c��D8h�c�"��x���UR��<�Q�-��{�[J(%m&�T�;Ҁ�Y}Q��ӦT��v��j�DPL��2�Jm|(3���2
l���tP(4��En�N��� 3/1��zK[�o(���b�9���kW���A�Z5��-��
����p)�=�]"5ۉ�C�Ķs+���ޑ )�)5Ւ�7*���{��df�#]��<����
i*F�@/-mf�'imƯ���ߔ��;b���1�.���Ũa�P͖������gBL!�h�rʬwU��=�#�>-Ƥ��|�*�D�N����[me�[3���I�%�p�������`�gp.���Q�$�f��IFf�A����`j?7������#W��J�L9:���YY$5T���2���A#�N�ݡ�+�{v��Y~�[���`g;�Q� 	��VN`��!k�8a�����;��oI�o4��΀��j���!��.�kM �5�>�<*:�N=Ԙw�t��=g+�x��)}j0��j��I�y����s&i����p�≶����*�<W�ƈ�%��)�̣0Wqz_A#�9�5�Ӊ�fG%�J�y�:TUF*��_q�b�T�d���ARÚ�{r'[��I��\{�ް��CG��EXxm��mw�G�A��W�73P��i|�$�,��A/<�T|�5�!���u�Ng�I_��Y2b%`�T�֫sҋT��o�Q�����[�4i�C�ÿ�K�?zM���"}gx�Ѭ�%$����|�m�PO��+v�KN�g�9?��iMX��!�SI�V�4I_�N��y]�)��S%ˊ��}���x��qMnf�.zWGn<�*��|���Y�.s���Ef�R_�[uA˺��]vh�	�L:;I�3}�������܈�B����F¡-��D�i��"�a���D,�Hc�r,�K��6ȡn������{�~E2ta��H�$�X����顐H��6Lk3JƬ�a?CC5�T�]�ai��r��c�4��Z|�����K��Dz�aH�R��f�Y%�O=�ޠ�Д�%�u�K�o];�Y�����TTTl��"�X�o�Oo��p(�lF��Lh&��~�w):��ƪ�)�%���:M�8��,��X��6ς]�����j��m$^��Jn"b��b`��߹�����ynnaeK�a{���%4ƴ}P⯒���F0�n �V>�Luޚ����H1��zk��"״�(ޱ�+��ɰ� �d��k�WYU]�����W�i=��Ӕ�~ʖf�[��a�����^�2b�.[��SŜ�W�k~��UF�T�{2~q��W_���Q�T4�J�H�N��&�7>f0
�	Dx�1��Tn'ؐ����M Dâ�B\�6�4�TM/7��"x��z�U��8@lA�\�i��)4���guHN:/m�w�z4���7�"J���0^��k���p�c�E�N�K�?��u�T2Ok�]���%oӐ�������Y�ѢCB�?��
��",n^�^2�,��x/;k������p���.م��^�ݭ|�L����F��
�\Z��M�I�EO�	�-��n5rcxCe2��
F-��S6����&����%m��~�Ώsv�n���兲ި^jh����	��x���/:�2S�&���lg�ұ��'�9���)���&�@*eAGs��>��܋�b'x�c���mK��h�*��h��+�y^2���v��(���ua���j��_���6��y�&J-\g���a��������a��~e��{��k��Q�b���