XlxV37EB    93b8    1687x��=�Sۺ���Wh8w	Mh,'!�ig(M������1�O��g;ޜ��ݕd[�叄���-qSGҮvW+iw%���F�v�m���ܻv�_ϭ�w����	��o��k�t�p7k=�`@h��{�鿦���;8�$��0����;�͓�){�(�@�H���e�n�n�N�6��_�W @���S���E�ҝ��c��<������$pB'xpf,g���ܹ�Y��qLC�� ğN��� ��ӱ0�ځ����Ӥe���A�d�ܸ��e���ȝ3_���gcJHn�@+��{s���~1w�������I�ȍu�Ο�h�!�I,�h0�j���6(:]Fw~�����Ü?�0�cF&KM�t�6=jØ`��L9�0"��Ȼ���N�m�,ȣ3#n�[I�2��eB:�B$�e��""�sM��oyu�Ƚ���?�h:>�|6�*+�`��Z��I�)��F1׳�z�O7��GI.h�G��M������!| ��na��@IQE���l����$�z�<<&�������@�s��V�������o:s~��{�M����2hzD �-)���9�k��r�������w}hF�
9���2� aF�ro�w ���c���B8{��#
p�g��׮gA7q�y��ο� �3�� �|]��<��4 8�M�p�aɪ6�ݷ�h?�0z_ϝ2`$��e���|�<9�$�o�G��;�I�}��
n������ƨy��T�"��?p����b��ƂT��8s\��+���2�$g���x��,�k�ǧ�����V�H��v�Щ�d|>N&�6,|��;�th>����᧋�����h��o}������G���{X��Ó�S�� �fӹ��S��w��\�i ��ܥ�:�	+�#�dy��wv�x���{�<2shD�s�yl��⇬;��۸l]�N1�O��K�]0�P��5C�2��qF�� Xe�!�bn�طp�X�Y�c3i���R����>���M��2 =��x���a�MĆ*~�'1�3�f8p���'�V��1�ܹT��������K����̐����8�sx1�p�qt~�b́��l�\��丸��7�+4��/����ۤo4�����$�}���H�����#�)��:�VjU]	�P�h�E[���1[]���Ӈ�!|�9���a��.�.�]]v���J�Z>���t��;b�e�h��]�6r�L#ϛe�˻�{+����Z�}�nA��F�E)cT�a� �t���n����@�|��Ohd����/B��o�$t=�3P0��a��y΁y|�y�^�c��^�C���^�t�@_�>A:Y��p9�
���h��}��2���86�x55b��ޡ\��H۲�G�� 8R�|��y$�B.	��O�.�'�L��W�[��2��l��
m[h F�L��ν���̲�G�b�ykߙ�ؾ������N�g�Έ�1W�n�2��c�3�aݗ��K��8�}7}��O{/K◳:D�_��wO`-�����%�����Y�������V� ��9v5v�l�@LFy��/K�5u<�V��=}��>�hL�x�N��U7�qTو&]�٧/>=��Ov,�G-�l�Zl�8e�f�I�dj��J�ԤJ�'�{�����ݡ�Su_<�uZ���A���"��F$�B1v	����nze�W��&Հ���U�-��{=�L!	g2���x.q ��_��_��*v�����Q��]�DWq�(�=e�R;�zY17]���,Խ������Aϣ�^Y�s�G����G���۷!J�j��������\S:U�CfԴ�@�����;,bn��:��v�^���5�@Gs��]niW{/�����.�v����\��֘ܕ6w�ѝ��TB]��E����ڻ�z*�/	ےNK�T��0��l]Ӭ2:O�D�mսC���^�+狤n����,��%�Nk���O���Ef�-*�mf�����X��`�_��vĿ��~�����m���F��W7V�����밉hu׍��>�o����^X�^JO湭}��Rڦ�6�?F�?F�?F[5��6�mp�C�̴�Ez��.z��ϴ��j��E�����6�G0�m�	z�[�Yۍ�hx!�r���y.��6�q��#�Zq,��*�����^�w߶��	�Fd�G�m�������ضK��n#`�X#�GW�ȷ�"�
�+�2n���o�׍�K�@n��I�<�H�z(�B��r#~�bnOvpci�o�����f�#i�@bg¶��l��b���#��߁>p�@\�D�1���P)g��R�����Y}%�'g��2]%�P�Rd�JΑ�c��ʒ8R�dQ*BC�q��)�����A{j�,��)KD�!KD��HDmMC������P�ڠTQ����R�j�RY*f�,U(T�**��P���B12(e�P�]�,��4���j�R1U��/��"{?�N���iO?���79��&|H�C���=���A�	~4��R� %c�f��N�1������S3p�O��[�w�+p٣&q6@*%y=��Q\OR>sb]�P�6�����D��I���j�huMT[��j��׃&y%�QȠ���Օ�M���-
/~�f�s.��9�+��@u)�x�'_��T|"1�6�F�s�x��/q3���j���H���+C'�5�0	��W�L�Fb���G %sB�Mn{�Z����/m�}�.O��2i�^ӓ�Y*� �ǩ]W�yU	�)+5]�|{�끶���9ZM\e}pM�E�-���i$M�Y�1��J�*�Cɉ�{�����b)�`H�4�2j�7�2�:	��MM���e%؍g�F���d�ao�^�����X N��O�6�����l��|�;8��>x�ǱقS��YH,b�f�)~p���#ׯ)>��KoʟE�߭ �;��9%�l����2Z��`�H"����[}��׾������ٲ�[v�v�,H�7Dw�f
�HW�e2��r�G*�l�CA̼����R�=�Bv�!�S��~V��!�!�u�1�,��ħ���ýR�1!��K�,��:�T���ȍ��HD���j�a[K�C�(8�bm�6OV����Akt�|�]���NRG_͵�� ��v��]�w���z��r��4ֆ�+��F�"$�j�rc��xwS�,��Z��DNU�B�zg��x��g!�5����.��J ���n��֐T�8����l�q�3�ˌ?:򊟐Ѻd�k�8�X䖖�i�!0FjW�ʂdk���j�\�,E1�y27���~�N�U�m�{M�4e�\h5�Iu/�1���OT���:����z@]�D/�&�\٫u}�F�+�YW���Sp��hyg�PL+���s�V�i~vX��������4?G�Fb��uɬ9Ov��)�#�C�#�b���!vC
��U��/qd{�Y�F����u��	t�E"���D�J��B��P�z�>�v��nzL���ͬ\�k�̏��o3�o'�'e��[�d��Z(e�v^=we��V������Ȱ�_-j���W<��7�rU�� ����S#�d���N�o����j4�|y�H����A��u��+��C������e�����F@��
��
��P@=?E|�����c9�x���M�|�Q��8m��f\�F�W�F�~��,\iCU�|�\[��a�T��^��
��}V��]Pz���X��y�����9u��*W��'���Y��+��!0����� �m���f{�����9�6M֗�س�ԊU�f��κ.�j�珯�r���J`�I�����y�H{q��hKԭ��ש���ژ�l�3[ژ��m��6�eݪ�l̫�|\�&���|�F���E�b��18j�����J�2��U�J��J:k;GkC�	�t��=����,�����K��?#XBK~K~�݇Zȴ�Z0�4i����m=��O�N/�{Nw�'uK��U9�O-zH�)}�8~���UH@ɟ��𻵐I�`�rhCF�.�iz�S���/}�;���O�z�b�������#N��5�쭮�u'��IKE�$_R9�D���j�%�	�cMܒcMxd��l�ɗ����Ѩ���`Xx�I�aXx≈�{�F�?�����p��#'da;�m1��{	iZ4�b��E���0p�o���S�c��<���3���,����/N�)��Qn����Pc~������|�!
B=�F2����QFt��(�I�s��*1CPHX �����Ŋ0�7�~�v[}�o�y��c����5�A�v;�s�ƕ�� {�=��r�;����~������[�]ۍ�b0����k ��×�b���ki�f��J�eL4�fM�t��ņ���X��FvP�{[�(�00�ȞTq���s�X�8~#�����z���e�W�z��ǯC���Ѯ����kȃ池D%D.N��SMq����)�-.����e�[���*-.��t�ER8�����){�h�pR�n��@�b��"�K�h*O���S���U�]z{i: �1��p����!�{��O�*�5@#7P�YF������$տ6:1�d����T;�a��+*H�`����պ0�qd��cd;��l�t�Ϧ�Q c��ێ,\<$ME����(���L�&�/��R���@J�l�)�R�1��i�����2�L��Y��:�*)�FF4�Ѫ�P�GFi�(+(sa���Zm���vۻ����ڤ+s�[���*�j��
MmfD��rr:�"��7r�������Ɏ�������xR��\iG}��e�l���L-g�<�8=���^�7Qs��G9s��ݙ��!{�705fP4T���D���b�0~ސ�t�f�����6�������@���07��%ـ>��{0ٍ�'�dh��j9F�G/"S[^=�)f�2�����U�������p<�<>&����$O��Q9��-���_��������}�t�c��l'VԌ��z�I8���D�&��ŭ�^E��P�@/�����؉b�Ѷǣ��r����y���?�jt�{Z��<���cLq��8O/>OG�.��G�C�wV`�k�FI�O�<M.�/��w�CЪJ�S5�:{L��Lbw�3�$#N�I���$Ɍ��IR7N�%I�8��$���$�0N$I�8�(I:��N��ڳ��	�� 횧%��A����Cڌ�%!��i	 톧�<��
�����gI�-������-`��$Z¡,�vQ���Gg�ms'ߩ�OG^�����$s� ��w�eC:j��~A2a��޹se
~�9V��쌃�*�8���w�1�N�F#�Ι6�Rr��}j�6&��ߐ��^fmV�K$V�/%.u23��D��=�U'hlj��,�8l�!��������!c�Ow�77�|"8���YkV���7z"N���h�����v~���Ư��L��؄�4���fn�U����q.6w������kߟ;����z�S�O]|�Ÿ
��=�8�q����T�jě�Pc�S�8�I����9N�Ab�ü���؛;�mtj�т 8/���.g��B��QB%$�j���8=�5�ҚY	�T��P�\�B�r-���	�6:�i`(��'�(*�L/��4��Ӓ��4��z�(ӂ�!Mi?���C��&�D� �zE�r!��C����e�p�?{�N~�^�EB���H�