XlxV37EB    1607     670xڽXmo9�ί��r@!m�T�"�(U�Ҵ*I��T�̮V{������xX Չt����=��1��^�Z�E�äG"I"���+�Ql����4iΩ���q���q�����:ǽg�z�g�pNXO��k��۵�$j�@{�oH脄������V�
6:��S�#��ƪ������	�o�J��n�P�mz��v8��I;�I�֟���<ygS���kO ��e�dVI/�M�W/U"�HF�җ�΄WF��\��IЕ(��^&�}�r�HK���v�.����l�`���%�N&�{��&S���Ʋ1qj�FF�7����B{��T;s���GAs��di��X)g��8�!���}��\�L�.�ggrK �H�$�JP�n�
�Lk��6y���Cp��oO.c!"��M��,�K*}*��exc���i�h�F��ٗЁp-����l��8U�2�t0#�^�L��k!�\�e�����Gi�{��^���U�3�Dn*�BZ*�9V7��a�}r.�-�*�R�h�h5nc�:�K�����R*|�'��R'֥��9����ysi]��)"����4w�,QM8E�a�A#T�&�+i����h�2� ��4s��͐�2P��KR�ܱ�݈�f)B�+��E�o�w�����oOڻ�]��P�S�M^h�vV�E��~.�!j�_xŋC3 ����K��E+������֟��C���j&]��ط���!&�w*�Z�doa��Q�x�J[�q���/~A�Fe��^^������a�mƲ�&�v9�wS��~jlo�}bpd2峜+����j��À/��W5��X�4�1y��3��W8�Q`hu���tX�;eQ_�} �OŌO��s���so
� 15W�����6V��Q��\����
�8��s�_Q��ߏ�V�����a@��[V���U�.ւ�U�0`bf������Ln����Ӡ#ӣu	\:Ъ57���ۀ������\y�|q�/6�1R���ہb>3�0f*�i�㱕�c�9ň]��њ�\���brpkt;-д����̆ʊ>��xR�U\��S8,*|j�-A���p��zpaOȼ7[�����0r�VϳL�cRE�5<L��$O�?���zh3�9�Z2nfE��f~98=�]D����G��;?��{�H���H��`��_m�(5G��O�8t+D�ϸ�"l*(5Y����v��5˂�z�]�<���[$A�u;/��|�uZ�Խ�v�g�5xKȜB���[EZy3Ǭjl��c��6
ѣ|Z�^�d���Y�@B��V� %�(���5ΡY�w�ݞ/sƕ�W����O���g\�h�G'r0y����D��
�I�R�C6��:����]递������>/V�� v'C�^+ʞ�?�[ YL=즗�8g�Uo���_��wr�v�r���S� �VBp�>\��k��C��b�U����_�
J��o$�6V�NA.�"�p���DC���Gm�q(ee���vH�^�B��a ��k@#Ba~[
�� �����tWF���4ﷀ�A�+'+F �M2֊��rJ2�~�����`��M��1x��'��ڸ,Rb-�B&�vq;	��Rz��