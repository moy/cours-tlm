XlxV37EB    1e27     64fx��Yio�H�ίh%��А��cwa2WB+@fm2a�H��;�c��!d�?~��@|�	�M��"��^������r�U�R�L�S%Sn�Z�0��9��͑�<�.�w�����J��{����T>W?j���$� �DH��9(�__�]_ξ���r��u���q M�$��!$C�ro��P�>%�u�%�! �L,�s���Io��e�5eյ�7Gz�X`>��E�h8����ꖍ��K8+�~x�X�P��p.T0E��������gc_X��Fgl����E��ʳ�j<��Ȃ���jo:<}�T���#�ᬬie�L�\p��;r�7��oM�7���̓�T7[b�!_0���$�c�r�*������xٮoO�;D^�;�{�~�_�?�/���Bvc�dJ�/���?f����7͓��f q�=��C§ˏ|��[;�	c9ddj��K<�#S�Y��gυ��@\�ώ���t�=J�[�DI?s��sU|��4��U̮���Gg?��ܓȗ�d���tY��l���b�q���"�����!��p�����j4�� Ho�փ`�i��.�9, #ȜGy�@nf3&l+`16��,�K� �~�lFrkg�'� ���r+jд�v@?̯������M����s��#a�'B��v��>��c���ۦ�}�xj�n�T�Y��3ғ���f95��L|�s?�l�Q��0�籩�? GpX� UB��@�i�u߼��[�׎�X���7��\@*����di��0p��>�H���q-���0�7s�U=�|�1<^����1�d�NԤZź����7t�?���T9�x�*Rɧ�`B@D�qLpV��p�s7���V-ԍ�h�L u�QKQ�((��54��L�N�H�2��<ҫ)��$�J]c���<O+Ͱ�<�4C���f��<�4�u�G�M������b-"wFxG�n��\0�R0�,/�I���`|wp+z�`�.}�^���ߥq�~��e̵�B��hZ �^�4��b��aR�n�2'Sh����>bs�Ї�kc5<7�'�]Ϯrk������vQN�lf�݌�W��=9Z �19W�?$����^J�1UWK|�܀m�k�S�22�}XX�ݣ��Ɩ���r6[���	�N���^�ٖFzg!/QZzCc����P)Le$�v#�,����H���З�����m�UJ_C�.�_E*��[�n�b�7��j�B^sg�w�R�쥶���������е0Ƈ 5L_�a�S��VF%"�U=қ�h�� �����Zt�2�;�ݵ�Ε@w.�{-П(�Dd����n$���j���;�$>�Z/��+;4�ت!�~���(�;@����x�8�%�{��^b��(o�J�ִ�q�*	/���.���.�����ՙ�j�+�-�$�H��"mB��	-�(���Z$�E�^$�ER^$�o�/�`�{�{���������í���-LG�q�<́5�f4�G9#�B��A�:)�J�IR�b��m�	ID�<]Jk*@�1�H��X0�N����uRd�
�� Q�j]��zL�̬^(F,��ү��A���7�?�R/9k�� [�x�