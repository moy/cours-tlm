XlxV37EB    27ab     8bdxڵZ�O��޿��4�
� �r�a����kiY1w����m-ҤJ�RV���Ǐ$vM���0�y��w��qfw�7}�j ��z׍��}@�m�vPH��c�<^,gnk�����_,���!jv�~�OP�pᐡ�j�~ۆ=�Ҕ�x���eo_p��(#�C�����-<{k�
t,�B:�1�L=�Zh�;����yH0D|H�$����W�#>��Nb�	N�	#�)ZZ�6�S�$rB�`��`����5BlF�0���:3�YM
GJ�RwL����Q���%rJ#FB4�Kٶ�!cώT`j,�l&�b6�l�4��g� ��[G�%��nk�}����i�h�d'�d����%����:����� /xE��؋:��i��~3�r��yY� ���?�K����O�f�Y<��&��S\ ��-���$��:V�a�il1D=rɄ��E�mA�W>����8!3��r�O�OVLuJ|U�9q�v�����9�|L}P��[�(��5�]O�6�O�x����'Ca�sʺ=i�9>������#똹�D�G�6 FK(�� f���E g��G3m.YR��"��[\@��d֢9$Bc�^)���ł���&-E�N"���x�ͭ]>���a�N,4���7�~����O��z����ᩢ��q��74�����x;��k{��:�e�`��f���	����%���n�m,9��b�\�x�)I��E��s�V��C���d�6|RS�|ѹT/ߥ�r��򷑓8�]�x8�;��)k8���Q���K��ૻ�/{��=���:�LB �I5%���~r�:g�谫�G������w�|��z���"M
�����'{(ŀ������=��)Op8��k$�bn�K�B��{)H�0�yX�Y��(Ο�qx�)w�xU��%TPA���^�v%�eC2d�#�n��?c��S񊂬rte�C8�NkWĩ��:*^c��a����=�,���_X5�b�QC�~���س�n���{(XCS�{E�n�~Պ�N�}#h������hx����:@���qG^A���{1y��$v!_�����[ɾ=����W�����yp��˚B6���O/"2��9e\�V ������M�~dxbdJ�l�rF%�$�+|hI9I���D,�!���N�����I�H(�CBY�	e}�'���\��oq����>���(V�¯<Z��'v3��8��G�"�D�Q}�Ôl�k.��a6�F�8���*d���y���\��������7(�,�4�BP�{�o���\qE]>�X}�*�o����{��SĉQV~G�2A�+c��ɾ��P�
��R�W
-Yɴ��b7Ij-1�ü�M�}Ƭ��*!d�NTg�(��g�<9D��;��ܒ�4���e��~��5�	%Xn?�#�3gB"�x�0�J��L��~U��L/��qM�����L7,�N�_���m�0��K��&/��o�(���T ����^�W`��N��WA������}��r���ʳ��`K�?/�:)
5:�:���x,��	.�0	�%�ڹGצa���3�3��ZhK}:ƫ6\^���A�@��	��]�ٝ���S���SxךN�LbV5ƕ��W�~�O��~<:~�õ�����1Pn ��� ��� |����E������F�F� ��
�a8����'!��IuU�X'���഻�3���
i��ẗ& ��}9C��-�U��r%z��3ހwp���ozmSF��7�Y.��P��?�Q�j%����L�P��q��E�>,ln��2�U�
���7�0�:��냿�&�s��ycf����n:-���Z�����{iU������a��\`�1��DDI_-��h������lt|������	M�%�KZq��F���4��_�r��%m;𧣦�u�Y3����
)������臮^P��� c��vKI,�b��$����K���d1�F�$�O}e�O�&���M�J��U��wQ�f+�A�ZݤGI�����V}ǝ��U�V�d�pJ��b�V\�.>pjYAkk^�d��q�#Dw+��"�yz��ވ{8�2����R}���]E�wQֆ�ҡ�����c�u1+�ۊMj�˪@�&\^]i��ܿf�����>��;���P9�Ř(�Hy�$���)i�G?8C�M]nX��+MGe��sDn�:�}�q ���JY