XlxV37EB    2e38     9f5x��Zmo�8��_A����SR�N���p�����S�l�,1�.�$��I��wHJ"%S�ӳ�˝?$�f��>3C�xv6�o����H�?�޷���~`<�nwQ`+'>�>��i��VՏT��ijW����(��(2����1t��_��!��N����'�V��aB2����S!��~�:�-���{�9��.�
q��-��)�gT:�R�{�w38D�7F���T���U�$����	✬oo`I#�!��(~���Rc�a�,��.��8c��cL�K�?��Bk?4=B���~��e:�ǈ�v�v� ��3r�(�~$o̍��ޖ���E��K�;[�\�	E��3ݨ�d�Ʃ�5r)����z&e����3lg�.������H��`�)2 �]��{8t�:Q&�7N������ W[>��
��*c�6&�/#?��QW⳨R�J��C"
r�(g���� %�tkE��� 8v�}~n^�ͮ�R�w�	�p��&�SˋO˰�̲rq�0Q�9d6`F[$��I$1
|(I���g��ֱ0��/=H���U���F��
<�''~@� ��eFX-�-E��A���?�͊K��X��&в���\��_t�ӻ��7�/O'��
��������~;�b�p��c�vyqn��@���>�%�ڱB�`c{a��a2������W�hN���YxN�l�8��rc�B gc�5C��w3��d�!':�sj�P�AMs��yf���G�~� ���2F�k}|GS�U�w' �K�k�,>��Ԍy��1� �(I])17�m#�A���7^�H
���{�=�n!��}�1Պ�q��fP���]lz�B���[�z�ēQa���
#�G�a�b��#O"�I$S�?�M ��ON��P;qc�I �!�������0vI�kr�C�g�a�nla��M�>�R]a��h׎�4\V��C��g)0d�Q�ǉӞxz��?�?8Tg���T&�`�C�X���l�m8f6��ю�4�9~���Y��!�f��{��A�']5ˆ��,4F��<PR���3Y�a:#jeb6Y̢�R�:?e�_o�Hl�ms��\xt�.X[k*36����l�6��:�i9�S��J�~qUq�B���5��[�p5J�^,�w�8sZ���^�m��2CU���I�i�:5֥{��L�wR��?a�.$F�)kL���f�L�� 4��pb�\8���}=�iW�A.ɣ}�G}G�A0@��ݯ!Q~��_�0�I��	�����w�������ſCi�}�3���j��1�ު׌*��@(������2jj_��7��3�]k��ڬF�C9fr�j�?Ȧ���Sk�{Z=�]O�Ԓ'���2/�@:���K9Nk��.:��UEҪI�jR����S���5��ꢃ�5�g�4O��-�1?�B���c��H��97�5?���	z�'=P�1��.�ė�1�G��5�h�ߵ];��Z؎v�ȴ�2�
$b�@�#N6�N��5Wإ����Prv	�ۚ.�"[A���r���{�<��5�^�WaM���r� �F��Qlj�WW��F3��M�%GsHK~ᴃ�Qu��ƾ秊�g� I�\AJQP�!�{KcԻ�,�l�7�k��y�x�J����F3EmY�;�t�y�Lȟ)S`��O�(g"��
�:)S�����s����~�6z���Zz���~h ���	qG(�e���)2�X���q�J_i�_��|�a�1Z��'�EO��؍0����(ǈ�-4En,"7��-�F�ک����a]B^�������mZhx���I��	\�:�L�&g�k� �N��U�"C�� ���������-AP-�d���F�R�(�<ʞ`jT��"�I�+�A�%+*�i��'�W�*+�ŵ"}�u��۶�y���*���wނ~���T�B+�	?�����I�[W2&��0m���0ЋV����-�w2�%�7�r�I�-+�]�g��<�%���ekŒ#��}!A+�>�`ɿzv ���k�($��e/H�<xT15�{-�&��>�l(��u_ziƲ1]x3���-�>JG��v�����ɹI�$wbe_J
=���ޫ�)	:�I��M�'a��q���a�,~��>hc�r�PZz�z��o����p��j��4�i��A�zT4L���h���?�������{�{Y��nQ�/� e�N�Mu�*�&�/����Rï��k��;�Z-g�_��� $��dWz��e������fj��T�k-�����N�
�%�f׃ ��l���_m�H��l�@��0f|��$��}|���?���+H+
13!t�Q8��e�1���^>�reU�����߄��������sEş��'W����'L%��Fzu��x���ʭV+m�{٩(�Є�@`��AB�q��Ǌ����p�����Qx�������Ɓ��C�Q������k�