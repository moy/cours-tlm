XlxV37EB    4dcc    111exڵ\mo۸���_Atp��IM'�n����8B�Jv��/�b+�Ne�W��dq��!�JQ�r��,���C�pfH��������s��6Qx�;���;��k�ܟ<>l{�����A���C���I�����|�ĉ�N��iO�ut��E��T#&�n�1!{g�ùw_�1l���^��  �p�y�	��|/x�=؜�f���	�$rc7zt�'���H�1����=�dh�-H�͍b/rb�HO�}����&��I���'��%$y޻1q�-�;$"�a����Ks��\���5�n%�a�"��Z�JE��@��m�}N�!��<�Q1�>�� ����$��ϙ��Ӝ��`�4��<�}%Q��z�n����jt`><���ػ?>'��7���M������Q�Ǜ{����o��oOo�1G�L�0M!xY
�����QA9~l�/���ֽ�w�M����K�����d�l K�)��Kt7�6�(��@�)�6����T��+��pW�����&&��<W� p�[��C��mc���&Hދ�\ڭ��(�[j��ր8�ޑ��	A/U�yEk[��۸��@=���Z�g�lA�D��y��+]��n�qb��-
7n�mA���k�U�}�4�^$X��T���W����n����^�����8��ȉ���iڗ#0vw'[�ｍM駳�����Jx��:�_)s�མ���z��_�oi���G�?�$	a쉳݂݁	�'����W␟a�E�{�^�<���B0�[/�y19���Ȼ'Z���c�0�O)~�Ƿl�>��;�#�lO�,9G�K��
�~�'-��
IO�p.��k7+{f�쑾"��:���/��K�А��L�8���_���p������\�W�bn_/�	[P��=<���o�8���ݗ��z81���@��z��+����ւ����p5���,��ri�-�֙AC33}�ݯ�����Y�%��MmĂ�mA�U��g�.�	�k{�l�T ֥~�z)�XL��KA�����-�� ��5�L1�~��87��/R٨�F���dr��k��%�b��*^a�|h�֖�_!�M�x��>_��~8����|�G��k�Q^X�����T���p|�aW�yL��j����}����U���n-�I�C��
j �ցݴ:��FNq�&�?�Y��?nX�� Ws �|�X��~��͢ѿH?��kX9]d�Kj�y�'��a7�o�"�ҧs\9m�ե�x#�6�gg���0�� �,�[J���ԥU���G�	��T����)�"�p��Q4�*�.�W�05�u/���O��˴a���B~2�oA��� ��E�t/����4Ȣ)dĿbS&��f��AL}X[��s�� �P,�j['q�΋"������x��d܆�3���2O��<����@�����%���bS�2`@���C_0v�w����ޝ��Q`�F��-���Q?��V�L�@T�L-&�̊�t��8EW�g��P�Q�~��B(�d"�fJ9y�%�����bV��!;��Zr� ��5����~����h��/	m1ۻ���W��sA�o��7um�Q	l�
���N�a��R����?�*�Ԙ�C՘S��8��̼ԧ��i����`�l���~�t�t�,�g��'��� �=i�:)�lmtJ:��� �o3��R���0t͝�G�rh\4�P_�1-%,�Al*5���3~����Y���[wn�h�J5�J�x�
Ip�U�2f�Y,ǋIk�Q��8M�y8�h�	����h^I9^�*a������]�N�q��>�!RųԼWA:�0�EE���$����YU&7��8D����kS�vZ�E6=i��MOi��z� �A+��'yra������=/s�����C��~����@��T�H�~��o�i�Ģ�{�9�m%�m�)��Q�:?؂R0�TY�̫�2�%�q� :���욯^¼O)[�%��g\��\�i�7_�J%��X�b C���6�8�& �\�P]g&�p!H�%�έ����Nlk�0����i���v��1PM�qQ�[��ۺч��:%�$HϞ�R�3^|�����w#��GnIɟrɃ���w�����0��Iw��]�����@U��;�"�տ�� �Gd� h���h&,b�BV�T^�w6^�'���iO&��m�Tk��[�64�Z��'����M`��W�e2)�����nMP�i�G�!��1V#���qn�RD��+eT֏+UTҏ+�TT֏Ҁ�����A��+������J����T6�J�T:�!kC%�t<2H"��9��2��IC�U�7�4m�˟yb[�J�)�!��zK���i�������]��W���KfޣUvd��/�����9+\��F��=��MCMSC��LI�����9��IO%��fa*�i���IT����Oe�����L~%�L��1������n����������!o5�
�,o�2����"�*,q�
ݓ�nMU��YN.�`d�+P�M�������
S���y�@�<��ʮ`�ɇ�o�*�oTg��ܛ���J�<ȳ�7_�)L���Œ֕�%c��x*�㱀Nx*o���/����K2��oTWҭww���u)�9�6v1����x����|��1Ww\-s�)?��2��pbVg��1�=����Qoꛧu�D�?�mL���:y�k�3S�,T�����y$���'
��k�/q6�7c���Tˁ��糘� +*&�m�傠��*��SjCK}�|�ԧ��.�ˈ��(�@J��M�+�W�4{��R��;�V��]X����*�E�P��#�t,��}�.�i����D�T�TM/.�KS)�h�H>���Rq�~f��P'/p�8	Ȳ#ŏR�&g���R�Fr;�"�UR_����F`��hCk-�bm[T�-/qC�<��77~$�\yzz�Dh�	A��$o18~Լ���b�\�1X���jw��*W9�^�R�c����m�t�^*�m�nT셱6�5�n�}�n$��,�ir�?2���MC�'�בPk5��2Y�92����0k�� P%_yYSl�J�|dh��SP'�����3Y�|�6�ª��q�W��FҁJ�Uu뗡ϯ�9���hx�b9�.Y����	��%�\���}[�4���3,~��j��j��v8̇�x���ɤ�k��O�pe^k�0��4��i�	�f����M뙥�a�*�� ��h[�0��.��L����j��i_��Q�D��`����8���ej��x��Y4}���h���- ��(\�u�u����=�K5��q�y١��5R�״b]���L[)Lm�4�)�iFI^�L��J�D3*r�f��5�(�K���!�Ex(��z^�^+���|e.�A�j̅�+�ZIO(����U�-�6�`
�^��j��JL���~�f�]P9�y&B�T� �]*?;!?�S9����O~����Zb�Z�8[�7ڱ�Y+�8�?�˪�� bK���W�rDC�c��U��ݏb�'|>��b�TF�V;�ѩ���h���e1q�#E ����U�> ˟���e�ꆗ��2;��c�O'�bz��كd���W5�!dcX�VT�A����ov{|� r2��a�j[���ú+�{%��bZ�gh/�n���z����P޽�q�+n�)OɶK��g* X�bi�M.�}�k
U� �R�2!?���~t!�M.'����8����ƅl[YJ������o�}�*��?�oc7׺�8�,��LM.r��d� ��;.,�z�A�{���@W��#��	G����j ������,ǽ.=v^������1{s��\�7�W�z�zfkpJ��O���8O=e�_�o������F������h�C������Nt���-\o��y�8�o� a9p;[Y=�G�����[2�t�E�jd�\࿉�C�x1[��=�o�e�.�v�>d�!�>:ð�_��	����|��}�a6�Ì/x7Ż�֊�TgXve�Sv?��[�0���ٕ�O��T����������)��+�f�F�L|��o.��^�[Q:�t���K���;�膡M�?~��J�;E�0ڳ�݅;o&Ώ郿�>���D.x���jψ�V|~�� �,B�#��5�����į�`��-~���J��d�b�<�q��Δ� �z��p��d���ٿ!��b��߸��+:?��Ms�=זE��۪�����3R���$O��?k�F�hy'�Al`	]D��Z�?���