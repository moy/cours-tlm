XlxV37EB    1216     503x��W_o9�S��>�(����T��v�l��^,�k+�^y�N��o�e� KP�H燬c�of<��V�t��U���M��@����0b�1KH���Ӱ2�F�3\��|�_~jԡ�g��K��"����"���۫ճ];�|�Tb<ш��8+qo]Y h�x�y45����
x2�A1�%8@�%L�YXs7�Q�=q��tƚ�E�b�1�p%״0o��uj�:,	4������~s3�B6�[�2�)1LRؓ&J�J�'��4�g�`3���&`�l+�`Bg\,�y덌N�jg�=��L����9�p�¼�Z��*�qh����'O��˦S6��jT/��b�h�U��:10���T�C��SP�1���kCR�9�~C�#IE҄C��ȳ5**x:�P�x:��	��<ߟ/�6N��mNa������l��L��4÷��,Ţ��]���t��	f����&;j�YR�R�Rs��`�٘K�Aũ8b(�S�-`�c&���F3G��͂.��A`x�L`*-�K>9������c�����lK�Ґ8�[�Tj��@����񍴐�y�����4�fA�/F�MO�9�a�h9���8f:�	��U���������h�ܵ���BK�ά@�ҷ�����G���{s���楢$�XS����^�0Aܮ����4_�ԨW�Rޣ����J��ŚF3
��6����\C��;��]�Y���E�vT�W��6�.GFL��ؓ�����|bȭS�-X�C%CF��aXdd��fZ�3+���5q��tq�����7:'썆�j��A���$&��,�����M�	��:��I;,P�{�����v�|W��L\/#�bƙ���u����L�ހ���[~x�o�A�۾���@�p%��.%#��VG��G�����U���Z�5����M���>nB��B6GԱ���݇�T�Ak��<�r������1�<�+ȉ�?���K�Uf�/����q�, ��4�n�(b��0��Սxe�	ȏ�8I�q儬9�@.XmY���"�C�b���^�Z;�kU��`Y*P���*�z*L��6��k1�'C�8���a�{�?j��鲼@j�RM�>�Ѳ��32Y�PX�My�3O��ۚٙ�µR��O���ʆh^����n��e��JS�V�m����v�Y��Y	�	�l뼺#������܎��+v��5��*[~�l�;{L�.*UP�M��t�9�"�w��,I��f:?����6���Fۅ���#�