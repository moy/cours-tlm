XlxV37EB    1e66     82exڽY]o�}��x�ɍ�������4�5����}2h����I���5����eEv�^��Kdjf8gfx8d�݃>�nN��fB&����N���V��bQ/�A��2�^�_��_����-�|���=�OO݁.�H+��L��x!,�m�y˫���`�Zek-�۹>�P\�t�T�o0�q~JSp47\�x҃�b� O���B����XI˄4�i�i�-�����c�X�=���)�dV(	j���p�D��4�<�P<g/�	א��K�a��r��K播a�!7<�x�^�2�3��K�ə8U�J�k�rmr&-Xv�1.zi��C�V,I�$�kΗ2xv��g�:���R%bF���u�1	�D�s�+�/7K~�`j����eo���%׉��ׂ���c�!�E���|�������^�*���>b)���h3��}�C*��|LS1�'��LY���
&�2�m���G�⣲��t����g|f��\Y
�9�6��b"����+��0�Wɣ(�$A�1��ט�'��P ��Rf}�PD�9q�3Z=��3��ފk��T�D8tȺ]��%B#	��4�Y!
�L��|D�z��?^�>�^�0RYX���aB�v�K���|F0b&�
����(���6�����O�}�nҋTȦ)�e�Q�^�šq��%&��,�ؐ�޿��Ŧ�"Y�"2,,st!jN���k|?�r�C��EeŒ�����!��ct=D�%[�a���6(4;�pk�Qza�����,��}X�$K��.����չkɆM�sp7~��B��f�­����W1��d3B�-��a��?��	��||�e��z�A���)t�ﺃ�d�!�/~i	�-[�~��z>d�a��?a���9��6����D�K-����V�~����L�zQ�����T5��{�a�� ����Ϲ�Z��T���伢��%��|��Ʈ3��ßw7M�*-R��R�$rCÆ���zq�5��OUQ/���j9�K���݁"=��(f"�Çm��s,G�9�ֺj�[�$��I�<���^HV�Q�Q&Gye>A�Q�P٢�a�rn����l	.R�:2<��M=j�L5,h��j�ǭl�9���Y�u��QŚV�D��,�w������~;���T��Od~�֕���>����8�����Ϸ�?�*R1�x>�9�p}�����$UsO���U7�Q����{����o��B�E~����aH�l��=T�ӧ�epu6r�w�5�CJ��B�h�D?rnt].���}���ު̃	��W	0��J�	�:�6h�p߫����O�I]݁�!��F�/뢵O�h�"̈́i�s�_:H)�FS�-�95wji4U�G������%�F	��O�qlPw�&�Y�\�s씓]�B���\�P���C����g�^��!W��������U���8��ե��n6E�~�Pీ�N8�8���'�h�!���s�&}[�[{�1���)� �r)�%5>���b�ۦ�������v��o��?���2�������Z����+�������7�h9ը��k�:�j�8R3�8�J�N�Ϯ��.��0D5Z	�g!���w~�F���:ըQ>Bp~�v�����2�gN����?ퟎjsE�1W���?4�U@�� 5z�Ua��n��̛�P�g��v^�Z�j/�[:}��ƂW���\�{j�QW5�.��-l(��y�W-��--����D�0����9�p7e�c�</����!8M��߮��f��4���Lxj�h7]�u� 줼I���)��j��vJ4g�f�L�o*�Jk�#�v؆3f��$t����> fy�B���W�0�}F�WD���M�̝5$���*sW{�|H�j��re���#��C��}S�^�������.��|��G?j���]XP�N.�ܤ6�.%pt�_2���*���� p�8'�j�b��G��ѝa����
[,6˅7�'PU(�-(���F�rO� �	��	�[*����D���O��1G0�G ū"���"���]�QP�*�,+!��#��e>�oyퟩ�u�Z� �\�s