XlxV37EB    3f7c     a63x��Z�o�H��_�bV:� �6��`2Rd�I�@�@�;˘i���m�d��Uwۦ��p0�՜?�GWUׯ�^]�^?�S���o�Y-V/��T��Ym�p#UQZ0���HQ;����\Ow]��P�e�~+���˰gDs���X�^?��L=bx+���N�#l��O<'9O�����?{hLMj��P�2(���4gp�C\�ɬ�W�Q��rCMb��	t���FK�:���ԶBJ��E���5q�.�p�^w@�G�'ѧ&ab�w�=�)�t��-f���O��1�=g�]�#6H���c?�*+��v6�D��A��K�����l�#t��d!�q]i�!pṡ����CZW�ا�3�Y3�Gw�/�5�x��,�m������	2��ȥsK7�J{�'�U��6��3.��V��mF����^ʛg���e�t��ω�m�
�+�Db[A@3�D-8 �uI���&�=��A�C���ȋ'������3V�Ǒ�
|��g����T7s���ĸ�Kbr|�f��ș���w�W��v&���N�n)�%�f�(���l7 Fk7�~B��[�<���J|t�ی��e�Z�G\@#�dn�xx�M�r�H���%q�%�4�6��mA������p=ڥm17 �ѩ� �3�ݎ������}z������烧�c��NVbtk�"Nx� ��W?ث����%�{�p��f�sjh�[�4�!�E]���}t�+5{j�m��E�m����5b�D*ܢ=ުA�6<Qb+���^�K=?���:Rﯴ��×^X'aM�t�ӝ9T�'(a�k�d�҄n� .u��v��G�a�s�o�}T�l���T�jL�I4���~b�ɱ�G)� ���+���Ԛ�%�?��M!ö�K�
���UaSdWd��{��m��篟���_|F��Gm�9~��35 �{��x�=��V�7�,/�6�5��u�Ϙ���n8����h
��Xn/c,�j1�
��sً�{�t!:��UC7�a�|@=��2��Ed_'L&��+��k�F�!��ŋZC�F#��ä��b�Jm�kC��X�PA�}}����IR�F�ez�ι"�aT�� �kJ�l�h�:�˾��0'�␅w���+����pD�R�>�J)��:H��n.���vK�$���ܤs��`q���y��>l���R߽:hj�&�-F�<�/Wڡǰmy�Լ5���T�nV��a!rŧ�l��ನ��Z
r� Cx�1��P���QD/�A�qJi)2L��g�.y^���mrV�k����"D�<p�����+�*S�Ec�����_�b���<����C�.�P����~J=����qYQ�>����!t�rx��@��Wrg����'s�(�,�`c�ܑ;k��U3�i@�ëĽtC��q|s*�"�W�0�ewi �� h�"�Y��¥j@E��J��]�b� jי ��q�y r��×/@����'��}�����1�`�����6�6Y�'��R���!�w�ԶoJG�$\�)�\T��I�`�x�ŒA�һ�0�I��s�E��oz�O�mpW|��i���WU�n�!x�脛5�{b-C��Z�+�T����}A_�(s�V��`�<ȲvQ��s	��j}`4u���"��x[���,h�<#q�?�vߵ�'�q�ޣ
J�,�]D���q�p�T�~//8�`���0t����
����{�_�ڍR��hX���8.�{�7!�າЗ��y(�q��,}_��\Hf����)�����տe�
�
�qJFE���p�*�`
�('�9Ddщ��Dl����RAb�-9�Z�X��V�X7-J��B&�	���.�O���e1�&���̔%�W��T8�*=!(�a��QZN؅?5+�&B�
y��/�Y4��H�W2
@.ޕ)ż��L.
N��OKa%Q �����I	����O�~L��D�H��r�e�^�/n���O�biV+��^=yUO�J��	>,�5S�&(~�;dbMԚS7���A$f?9p�; nJ�� ��rP�!��&0x���%ҧ���T�yt,u+2��WdukR��F�Y�i	{�!�	q�*��%A����b\���=pQ{�,{��#�$��b�,@R��� $e�,¡lL�D�����߭���Zݰ'=�{ҳDOz��{R�������$��H���+�z`�X�dv�2�������������}4mR�]H����7�p�'~�Y��ǻ\�r�y�x�W� �u�G�G�o�Տ��+���B�-1J�o��;��Wsg����2�����r�34-2-A������=p>s3�9Ҝf\���EI�(����D�ˌ�pl/����S���C���\�[�Bک[�}a���$y$t��dE��|��SsGW�L�f�$���$'a�=�j�9�km]e��_��O����7���)�����29[��ިL�yV&;d��O.0�<Dr�� F��˒�ը��?�qa�W��Z���<�o�D{r�fQ{4�ڣ����p��?&��?��� ���m��qqZH��oX��������v�qx;w���������o��#�-���u�