XlxV37EB    1755     5b0x��W�o�H��>@.PC�<�6%$��/�;������ƶ�kU����5f�W�\��~��;�����̺V�;7�W]����A��T{���;Ƿ!�G�Oq��>��'3h�д������&XM��'�:�D�$!\@wûC����{.7s�Ρ4L,��M���H9=�Uix�:�s� @'���'�,`���Ы�n@;@�4�|F��Zy͖��АL����z�H��',
s�5�E��9M<�b�/�c�1��ԇ&����1�2� Uo����OUM��@��O��v*&_��'�\���w�^��e�f�֬OR���D,��ސ)�X��L�1
;���Q�'H�8$Abö�|�����c?@���G�D�\�͎��G��*]�7�%�0RR�p/+����3oT�;�K����Gb!�ELw{>x��Hl��`K)�t.�+{K̒�8/�ӱ�8��y�t�B�����(���0f1�HNN�X���,
j����|.'�c/��e��f�}`�Qj�c�
�L� �G�R�����c+k>�1������#
ḛ��g�/���#���c�=�PC�<�$�9�����m���SG�,�Bd'�]�����{渟�~]��t�޼U�6�/��v��D=��A4f��h�~�� h�����( ?�;��Z�K4p�}]���^$ݴ�煝~[��6x��M5X?g�w�}�����țo�\�5&2.].;daDv�Pڻ��r�e����%?��'б�&	R$Q�������C ��=6�F�:������{��څ��ӄyȵ~�rEL(��n;c
�{��d�LѦ�w��o�}�-pYR*�*%��y{�v��_]��v�1|�e��V&+�����@v�/��{Ѿv�ԄZJ��ig�5�eӇ��U%Z5[턒��&ۓ�_�>0Ó|�+�<�.�U���k��%�<X9�O5�V��}kz��(���E��b2}ؒ�ô����	��Y�����6�%�+X�O"�h�ʃƯ?���jK��F������,] ΍3@؈�,ز��e�*gY*����L����iƕ�Ε����)[t���k�\��!�@���E��P��s�UXS�iǚ棹V�'
��֓&M��ɹ}���>B�l_̂����Q�D�\voܫ��;��O2&CT�(��S�İ����F��~�b�Pc@���(]R��eW��*0���YޤNJ���A�P[n桲�\(j�;��bm�im��ZUF1V:�ۃ����HU��1AȥN��1�\�6Wd��/gД�#��6,�6�}5VE��[�B��`�W#�o��?�K�SÐ�,,�7��rN�@�)��Pm���y� ����Ae����L-ɍ��b�&��^�9c����o��s�U[3k��Ƭ���Za8:׈��ᛪ