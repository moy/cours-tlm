XlxV37EB    20da     800xڵYmo�8�ίѕ*�M�Na�R��R߶�U��)2�VC�%������!�!I���[������ػ�7�__\v�^��^��>�A}��;�dpw:uG��/&~k��m�:�b�_�m���ёcC�I���C�u��aӝ2�
���8�9��/$�&�S��c
[�X̽��V<% 8�f˘�'X����Co��A ��X�xA�}9�;&m#$=АL���a3e��O',
3)X���E��9M���x6ܟ�:��&`� ��T3����ocu�eV9js�¥nÌ�9�Dq�<G1	�ȟ,�Q�t�m�5�����=�H��X��U �d�5��p��.DIFa�d�"g
A�	�$H(z�nX�P^y�� ���zK�q}��Y}�y����ߣ=%��%ǏiHc�UA����`s,X���|9��+>�v5$R)�0%Hk!���r��)�YR���q��(�"��q^4��`*1T8Jࢩ������<�t�k��P�@ǘp
ɷbR��B����8��V���T����P� z�h�gs��,���|�`�E�աG��nA�of>�rh#�\/�O�~6��G�i�#�&	}K#�q{ws���΢P����N�
t��{=��o}������oN���b/���v;5,�i?�Dc湶}|�O����^1/�F����Cײ\���������P��R��z��M\}N%�@��"�|�$V�xg��g�+bI��Q4j"�g�%�]t������N�����w:�ȣJG��S{��Vrw8#�%<�Ú\]m��{��Y�����zL��Ӊ ��]5�H�rpE%a�&�Rh�O'�r�{�(nX�#��J��<p���n��M�B����w�L�w/�]�|��9����29��$��r݇u�P9q]����I�9-�[�҇¤�N���m�U���Uf.�W�b�(,9�1�Gs܀Gѫ+�{t�`x�g5��9_�H�-T�c�{�U�%�&�(����O=I�U�Lʒ�B�8�8b���KG�G�5"���:%A�aGߗ�#�{�.J�%�k�;P�RMn�t�+�Y=��f�ϙ�ґb׭Tzo5hW�=���鬃����������s e#�+/�4�"�r��p惽��E�(���R��6F��0VPa{��p<�x}$������|>��<��V�>��������̕��2���hcH�1n�'߲��U�_|�fB�x�u��h��0�we~��І6a"cq��3����2�^A����Z�N!Jn�j�@e����s�(F���r�9I��9���=��J�U'/���C�Z�Q����/D������M�h��#���|렎u��כ��v�%m�p'T߇�:�bx�Ε Gj-/����^&4�0���$oK�H��P],.3"$T�і�_Otո3����CČ�+6�����Ԩ���e�e��?�C� � ��81`g?��&a�-aK	[[�$���C�0�
��B*��v�����U����� a:X�٩ޡ̌.��A1�j���v��{S��Ul�_���b��icX�w�!$ϻV�zuH[@��b#��Y޺7[��ӷ٩�e;E>�QO\�=�Cy����%y~Ju��nc���
�A�=z� �%���A�tGFI��>h�L��OH���~�>����ͨ�)��ff7ڇM���Jh:����M��B6���#�5Z���9	�%fk�,:!�,����;�zX�:��������euF97w<dC�F�ETZ�5��|�ŭ����p%Ҧ�J�jds7��t���[��׃V[�W�ϧ-V&\vݠx�VܹΖiKb57Z'jCT~���m[�~�2c�jc4�tN4��O�M`s��
6/���=�l�g�w��1���M�i����EV�*?0 �����$;�[�&����h�Վ5(wk@�
������+�bW�o���4Xz�5:�8���!g5n[�Y�4����1.x�O��p�)����N�