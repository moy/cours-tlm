XlxV37EB    b086    1be6x��=kS�Ʋ��S�Tv���=)Ȧ����k�6�(����X>��B������=�p�I��!Y�t��zzz�1���>���!�g�����@�m8�G�����y�����,xD�wPww����vߣ��~go���Q�GY�OK�������1��xQ$��Q6�O�xZ����ĭjo�O��Yrw_��d�,�4\L�!;Bo>G!GY���c<{Gj�t�5�8�ǋ�!�/� �	��-��$]T ��nw7"+��,YU�i2���y�G��x��5h�H
-f0wI^ 9J�8�1�q��k�ZU�=譊�4�S���,Z��_`F��y�v�#�/;;�{;�0�q��E���d�k(���N���f�]���ݦ����2Yܡ��y?74�q�����o�1��bT��t<BI���F�%���3�����'�E8O��+M�YD��G,�E�_-X4-��a��'w�h��#���p�YaM�����bM�_7�p�<~W����M�3x>�`�0����ŋ8K�.T���h+�h�&X��y�G>�r10A�1z�@�.b���
Z�o��܊7]e,��"��M�����h�(��>��d����sKAc�G�@�}'5�Z`Ⱥ5�|3]oT� �w3�]ȸ���^�[`�H�#JoQ�*��-S85���6��i�\��� F��Y�-�GvN��������r���i���,��y�Q�n\�����X^�e��l �("؝ݠ*�O���p�%�y����_��~qQ�1On�({FI��Aȿ��Ōʧ�����]4�pXr:���)||�������,�{�N=�oM��+��`�x:�2:�/?�TT�$�ب���?��v��<��]P
4R��z�^8�>@���*8p�b��-ߣ�O��>�>�I���������ce[�,�{��Q�¬����-#A�;J"/2|x(��&>���颹��c�"���9�#P_�q<��0n��/��z=	{GG#�y��.��,�:��.&��3�w9��l2�./&V��Hy�~����# ��5��&M�1� ~20�d�3��1���9c] �����hp$����$;R�G���ռ%���>F�Q6�ep��E��' u���#<�t6y|q�!GZ�=�� ��YD���C��k�.��I��h<�D+��U��:�[^Ft� m�t��|�(?V(G������wx28�j<�[9��'ó_�J7H�6#G�����C�̿V����,�Q�x5�Zy~^��>Z-��j+�f�X7G����h���f�r�Q|�x��1Ͷv1���/w
��m����P�ؤ��X+���Ng�4f�3|x#z��ڎ�w>���/�X�׈,�_�jA���x<�#�a����k�
,��@�1��փ�
����x:<N3>�NM�n(^�!0��p��x�B`�:���1�����/��Qt��U��F�]�[��¬f�p*5(�X�T�������F��h~K$�����\����|�d2��#�iŖX�`˺���xF)A�p�>c�U�2�0�g!����q�z�;\�"Ҩ|�rJ5��<ZS&�#<!���l�O�1�?�w���F�a�����|��"�h��10�o�b榃�����2�cH��g�P�-<]=���J����c���heH�hf�+�{��ض?U �ڴ��c��xhsa;'���!ә+���=-�(V'1L{	`��aԡ/�=�=���(.���D����hn�Txf���@�=ϡ���OX��x�V�E��o��o2�ep��1��4;��$���@�&(z���	�mxQ�Y�p(�{�8*O��̃uq����1(��'ؐfi&���I�xL��x4�g.(i�+U�5����)���}�H�E�,Ҡv�t���+'������γ�s�I7Ų�ٱKW�� �j�b{LH��.W���e��oN�Nu��z��3|߬����w\�Kʀ�q\L�-��ȟ�}r��z_٦	z��f�����q[�'Y4�,�%Y��v�:�T}�Md��`��KizMm����	:I_s�wR�M��7�;��Y�Y�f�[jw��;=?C+X����l�p�<�M!)�Qt��28�@5�J��G�"�
p�b-�~(_\J��66~Or������S��������'@荅M��^�1�r�l�a��)�k��pO�c�����u9 *�F����qB�P��dX/�B�����T���3@<V/>p� ��X�A����Ñ��f����)��!,��hVf�J�D��`��v%��
�*$�p�m�M�/O&jO:e#�ҟ������vGM��,��J?��9�z�D~�M�����օ����<�&@���Fk��t��nt����@Hk#z�җ�ʹ}�����)�4�A�bs��u���xu����@H�ߚ�V4P]ٺ! i��2<��'矇�a��>�ݣ0~��k��� ��}A@W
P�{������ e�/ؠ���?�i�4$�g�ɥ�:�aGU�$�{����ѥ#���C+�{���bq{Y����fq��A7)�}L-aZ!��a�������*0zS�Q wHh.Q!=jj��z�6�9k(�Y��SM12�u�|zy�+���Eew�N�TW]hּ�`+t���Z{qC!�t�d��Zn�&$��z���\`�J�A���	W��A$^ȉ/��鄖��?��me�ˀ�����O"6��܅O;՚{Esuə9������b��3���-���v�uV��A`yjWP&E�8n9�n
<!@�݁;�q�O������9JJf������f�Ppu��-���j��x�^AA�Wq����RI+��y!8mm���'<�@ݡ�#�-��O��]�Zf�bqT��4�ڇ��)���8��q�S�� (�Wնhb���-㧄�S��r�12�Ɩ7c�L/��6��a��Y+o�05;B��nk���j��	ʷ#r�����[Rڗ^�L��j	�����[��/7�!�.TRd��
"�7F�a����<�x�I$z��������1���_�}���(F��� )�� �oQ�k@�%*��D#�S5Q���ߖ8��<�>�6xݶx�>��߹^�f��M˶Z+��a,g�hN�xNQ"��|�*s�䲍����Ơ0ctk��[��2ķ�mW��fUE�ӡ��7?�|T'K��/����B<��2P�Z�XڵT����iо��_L��q�hA<m��IҊ�Nl� 5�v�T��mp��h+I%��
��4{�tj`�7��m�9
�1)F3wS�16����q�zO"@���D(-�v9 \�\W;g��AR���G*(^��"Dr[(�`-����2���*��|���0�y�M���R���~��u Cր�((��v���%��Z'rցj�-�Q���;;�I�3M?)��р�K�>����%��I�=�_D�;�ͭO	��ۖ�p�YW�TԒVv|�CZY$��ѴP��x�D��.��&�W�a��3J=� Q���N��M0�M13pFs�*=�6�2������L}���_�$�^By��d���u�X�N2ٽ����/�OTx��d�bzy��_&�.!�&�R	m��	}3
}s
}�
}�|S�|��|��� ����AvH1��f��e��J��}?�w��KؙZ7���˩:	9e��,����b����78x_Xb7�j��zy�hN��m$�sm�!r�o��j�
髦j�@�Ժ�循.P5�U���jO~ռ�-4W![�9��y��=��W�~�Rr�i!t�J/3��ݰ=��f�,p����˶�ȷ�MH�1K}L�k�!Z\�`���L(� ��TK���p��rU2��@\kv�6s4H�Ç�'��aS���^�Ӌ2��^H�5π�Uk��JѰN.�%��Z�CN��I)�]qb^d��u<6���p�
,yPF�Zu�����f]ϟ��8^�-V���UP��,���2�8�+7����(𴓗��a�k�#��ѯ����i<g�MF!��zMc$��\E5-�+:*tPɗ*q��ML���&��f��$�����6���c�l�6m�Iͱ�7�cW��fM�r�ö��B��!yG�U?K�A�j��R������ί�Z��{ts���-�Rc�?��6U��v��D���OŲ��HAxL���x���gZ>��w��F�<��0e5��N:��2%�W���>dϠ�����@��P8;�-Hjf! �a[�K@و,��IA2�+G�Iab�c-&�k�R�*�n-��BF0��%�I�JNó4���ݗ�`?��`D��`2?�r�N��s��Rk�,_��T
�)/[U=����-���O?�?!��hX�6ܗ		�5@I���k?cS`0:�f4U7C��k?O�qIS�o]�������'����}Pɯ��ʔ�k=Y
�U��a`kS���,*��+p��N�+Q�A��� ����g��Y�UvlP۶|���S����-T鍍
i[t`�Wٿ�9�KH��$�!���8V]��8�n#�J��H�U�+"EI �$Ĳ�恣�A*lY`lY����`֗i���-h'˴T1BQ.Ld�2�(�YѤ�2�&��녮��%���UQK	l/��c� yI��"�LK�m��H|.E#�]���U~ ]UՒ�|��Z2q�y@����+R�C��{%���9%a�iC����Pe��-�.��P�Ɏ����H�'-����X4��}��bU�'-�JZUU�}�_L�B��
�D���
2��-�7�%Uv��}���*?��ΠP��T�vI��0D��Bޖ��!�JojM�k'�]�lط��$k���BUP��	�P��jb�qe��ė#c��r�*�-cS �T.r��N g�r���5���-j�����;|�/s��\�ꤜZ
�����˷�l�ĝ�mQ��r&*�׼ p@�n��c��� �ڪC]��kGN�r����N�[kR ��굚[IDR�X��/�`���/��M�*)he!���=�cP/vH'%�t�`ӁC�!�8#�,��pd��̟וdfq�B�̠�(:�z�Ҥ~4�h���riP�ن��A���S�4��0��ǠF�5$�0ܽ�א2�G�K��F\�.��1��b �K3���6w^�e�R��������jk�xCN^b�t-�R���P�}`9J6�$D(?�Y9�/���fҺ��H�S
X�L�^c�5��k�n}�V�rI[�5꒶N֖�� o�uG�SM�������|�&�9�)8G!g��mX5 ��b��nT9�<�������k��0-r�04!=t�J�������E(V�7�ꎗ�����"�����@ ��.`�ל<� ��?i�Ǳ�A��畿j�Q���.��-��GY�l�F@y����m,8LN+���Ϗ�gP�Y1����2j"�'��.^��mP۪x?mt;�e�ڒNTf	1n�jNL����gK�@� g�w��S�-g������njH��WD�U$�`�	\93�"��
��O3�Vc_���bO�H�@xy������OI^�o��&'� 7���Tp��U����k���2�~�`Q���=����qV�5��Q��@�#�4Do�$'�����V���bz_�e��&@��#�����N�n�+*��^R���'�m��;�B�ѷ�Ћz���k�ۓ%šA�$%�+.�`��@IHw`��%!�:@�W��N�	�����p��	6O�)ͩ�P���)#��F
j��t���иQ��(�h���%�� ���J����خ�QU��c��2��R:,G�N#�y�
�:����#BXf�|�Q*����� tv���e�Dp�O���5|��Ϡ���\Q�.�S�̑�^
K��"�:(�K�,����*�T��y����|��M��n���R�-
�t
���m�贁T_4�1x1U%Ʊ�=FLM畡�t�K��.FH�ٯ~8l�u�t�2�����-���N��:y���d�7���e���Bz��a�w+�	��Zû��oOOx�	�W��2d�B������5>�!����&�:җyHC�ې[��B��⹜m��o�E���&�1����������Q�PSE�C��G������Mcx��R����X���N7��=@J�����SLU<|���ω����^�����L�$��:����pG���%5�-Z����ە�*;D~���Q�Ś�Ɔ@㦖E�Ӏ��.��"�Vc�Uε��� �?��'�흗5���Ԡ���<|Kʡ�-���%W���76<�CZ�ti��,C���n"��:��x�J�n~��������}�,$w�����JZ�ɗ3�^Z����^jD��6J���#��%�=lP��NƧ���ٸ�G�RK�ڣ�!H��	�S�'�aT*�q?Sd4j'��f"�pJ��I��g4;�!����P&���;��Z�.C�Y{�La�yi�ڋ�l��� ��l��Q���F�P㛿D��^��5<o�w�P����Ui`O�+s��­[~��$&�8�+�I��:W��t�����-<��^xx9>9��^����;�*7��ó�HET6?k���{�����a_��i�<�"��PZ`C���uA4������=�;���@l�����#��&�$��s7����I^G��J�o�
]�I8Y�����}j����]�Q���:MH�1���V(��W�����+Q����;
��P+Ԕ�Z���+�(��(�y�u7͓`;|�wd��].l9�Z����T�/[!�2�f)�<[!�Z�R3Ӽ��F|�V��d�2]�Gl�WRV�_�-Q��ڑ�ٓεl��)\���%=�u\>MUY�O�V!	ҍs �t��s�~�5���5����t*��m�j���>��������K�