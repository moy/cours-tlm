XlxV37EB    1776     768xڽX�o7��_�*�ȀB�Ni+M4U���*I�n���3`��o���i��׾�#����݇�~?���t:�4::�Y6�[Z3I����i{E�n��z������3��>�����9a=]~���yx���C��^�5	����B�Rae#����=�>����V��9l�\�tM��L�/m�K�d���tҮdڥݧ��A�����r��O��^(�(�&�Jza�m~;S�D�D�-����^Mf�i�`+U�[5-�L9��+t*-e*��I�Y�����\�5M%N��{�%&W���Ʋ3If FFgk��
�=yC~!��tw�C��V"S��I1�R.�2�Q~���{�}��^�IՌcv���DRɅ��"V���gk�LkP��!}�B'��ak���\�JD��*=���
��BJ��M�^ӥ񮏀�
�K�H��rG�Rm�c��y	?��y�l�b�Z�yn�����(�xm<�o\`����'����T:�
�ݛ?�B�ɕ���]r�*�"M1j���u��.��8�<�2�#N8��x/w�[	{��ѷ�֕��EIM���Cd���&/B�1i¾��V���?Y%m\֢J^j�m<-�J2�9eHAY�C�%�m�p��q�ЬEhw�QV~Oz����{��M�.w���(�L�F�]��h�D!�ת�{���ϣ�:4C&�A1aiY�A�h%W<x\��C��o�8�*n*���u�����y�2��R*����.�*g��!�����u�e��^~q������"p��>�F��~�R�������a�+�J�M��o�0�=�E?��7���qY��h<c׃u�GA����s�ky�,��16�w���X�>4zŬ�i����яQ��rj�9�{���t��6R`X���T�}�	��&�Z=�>?�r��Sd�-ʐ)V��e+?�ZZ��%凓Ӛ�%آ����׹<�է��5I�CKກ!�y�W�=9s��Zf�_�B.��%f9�
(1c?�(�3˚`�r���@����!�亮���������4���6,0����C��5{��1G�R��y�)59����Iqx���YzHaO=-�y/Z���a�"s:���<�6A�i��i��O#�x����r<�-mn4� Q`�N���˷W��O��ɳG���~;|��"SS�"�.///���|:��\%�~���.&�E�!�{���f���t$5��X�-i@ paEֺh�
��#=�(�䘶�VPgl���5t�An�;,B ��1 �k�b�Wp�
�И��\��]mj����?$�����F�U�x��[��jz1�X ������uF&8Sk>K����:w�Q�:ɗ���4��������˘�R2�}�$�jռPx����|c�;�þ��2�YT�"����+F�ra(L�t���cp��ᚄ����Ϡ����԰�����T��@�B&���UM�X�^�fDU��D���Z�IL���sj&�������I�>޹J����#X$7�
��Ĳ�,=Y�d��	+���$p�`�j.8�!@+�S�>B#V��;57zSB�8�#�F� n(=�8|p�{�᜚��V�Nf�Q���k�`G� ��T}�����l��VY0t�d�&�P9R�Y��|C��p�.�V�W�Ju�� x��X��f�^����8����t0���DVȐ�����*����^���z�s����1�.��J�`��bU7�AT�������m�����f"D��f
FӭEt�n�?M�LF�������ˁ�������cgӘ�S�ύ�0HG@C���[�1�xD�}��q(wk+��]�8����|*l4�n<�/�6��O�ju� �Qq�E�~��~Z�iw��ת
C