XlxV37EB    3a29     a41x��Z�o�����b�[�	���t$J�,R_*t5s�VQ.�&MP�v���y؉���;R�fH����}�٦�x�O��@;�YM� ���9�Vw���4�7����A�QS�v��(��0���>,�N���6��c^��M�W�Q ��_<��.B�����ȳ��w]D!
p���Ж����:.��{�Ml����8�g9��D�����f�5Ƒ�ͬ`Fdɋ�O�װ~K;Z���ErW^܈�2��n���,��\����N��L�Y+�]���F6w�l�愑<v�˴?D Z����u�������W��ºw�9�
o�=24�n�ˎ�F����ܳܰ�d���US�����r C���>�2g��]���2�M�A���[2�{8p�2(��=��y�f����E���|���CB��0���;�"?D�UW�P���0�=p6������Y0��-	���p�,�K����#�ٵ5 ��:\zDr]N�{���������P����@��<@�-��b����s��f0ImNz���a�kG|���!�B�<�Ӊ���b��
1�-�m�x�F0���rp:��]���ȱ�̓?�^LF��旑���_Û���/�3��9�^�}:����s�65�}`�n��ʞ;v�O]�Ol��f�iZY|@_��W2�bM�E`��-�@k3�\ӿ�M�XzP��Z�̐r�W��"=
�
r�JZ)P�Bb:0���o�G�=E]�k��=Ǩ�"�Q���^,>�_=���.b��>:�NR:C=7昩=a�ڜ�@�Uf~L��%�=�V�����v���W	#���8�̖kZzE�������BS�0W؆�Tk�`q�lhu���#�e�r!���F昦Hed?����HERk�<�M�͂ ,�Pn6r,�5d3$h�bP�#L	�_�j�����G�/43���a:6�m��o�I!'�C�C��!�O��qY��+��X�������s�|0�g`�'z�;3s�D�ѽ����J�&�o��u�|[-ߒ�w��e�::���H �F���.+��?]-��&a��l<�]|������ͤ�V��:���b4w9n1�R��e�����
-��EW���-�R/Eoz� @�$�]��������j.2�7߆�Ih�����Z��8F�)񌶯q-CƉe$����%�)]eL'?Q+���_���t�>&�R�YG?ﰇj��{�v��:����t��&����S��4����>�8��JH�ڂ���bmN�͋�LW�u��؅�Ρf��/�4�+kL�Q�Q=y+�gd�mQ���$:�^��[ض��`�~vIj����\�_�c3���5Bc-h�Q\	� %�=�׈��"Js�a\�p�{��'�W�#��#���C����|4�����Ȟ����;����ܢU��g�hh$|܋:Wm6�u��q$O�+�8jn��&M��֧�{O!�D\����5�z�=�iWX�k)p�l9��ABB������sM�L�m�g�}���̊p��[�1f#�;�}�WIg�4��]����j��0|�����e�D��3�;D���H�j>hBt���de`�+w19a�����g@_�]a�����8U.Ͻ^O
+��Ԗ�^��Ki�\;ai�[ٓbZ�>Mm��\�i�{,OC������&�� �����%��NP[1�I���C�jѷN��@���tƏ�a�q�?N�m"׉A�rK�����p�|�B�(���i*DV�?/e��ȚF�Z&l[S�ķ��tR��"� +�J��[v�kM�K	I�9�W{�z)�&:V;%_iTb{o-R�\�tߘ�za�/��8��Ł��H㾨J�x�V4	t "���F��[�	�XZTS9�E��)9&{��$���$�OHR\b�7I��k%�m�lgQV�����MٴQB�,�)�8#l�:N�#iiM�WGYQ���crҫ��W+	�����%<���Œ��2�_Bf��T�j���G�%��I�sSj�X2�Nn��N���T:�!\[v�5�u�Qt�ِ%j�B���<��ء@c�%qꨜ j�C��QdvJ���������7sx�������1������_X^�x>�z>�|��3�n-U�5GEpk�&Z�q�P��%u]�U�6Q�[Ft�<g-��%LJ¤�t���\���T�2z�Q��si�������S9]CO�Ƭ��J��卷���[�����Z [�%{��?==�FǾpN�.�E=�/P;��mC���W�e�5�xHn�l��_E2�u%@b�@�	"9[�D�[R%/b���Ҕ�{VM�9R�)�.#D�k�r�ɽ)2��SN4���((&�'�=�m�F��D���H��<j�� �v�o;���l?�F���S���o�ڪ!#�|�2eH��'e��-2�����^�x�^�(��5#����ϐ9%���kF��߷���_�M����J$� Fr
`�>*O��(;0�n�~��"��7E�K����%�x�M���ZIz�)z�M#�e�E $��O�z����iF