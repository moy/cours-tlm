XlxV37EB    410b     a75x��[{o�J��O1�Wj�Bj���"M%B �Z�@*��jd��ن&���{�a{�Ĥ��{����9��sΜ瘶Zc��z����t�k���`>��>� �����n�����*��죪~�4�h�O�:�'���^���k��!����"N`/�\Z1��G� ]3s}(�
 ��_<k��Բ-繉t�<Eŀ�m#�G|�m�������Cl����c�H'�A�:��x��:�0ڪ��bС+⛞��a}���
��G*�9����%�۝+�!�ކ�Q�/�\Q���Zx��K׋U��g8t�w�\��c�RԖ���UJ;�<?@[�v�A�"ID��|N!���M��r8��YK��{K�Y�9���ˍ�.Z[���\2K��[ce9p$gKs��a0a�?�o-��;(��N=B��k~/p�i�7�ϭ����zl(L�*����p^b��8ĳ�2(���	��Ѐ���r`_��5)�|�xߗ���V�O� �<�Q'Gg~!��xlGp��3���r�b˰KEq�J��5��|�j^�'0�m�%1 ��nJ�kO�L'��6�m3���)�DZϢ����&Xo�v!)J8+^mN��I@H�|�4�Z`Ν���h�A?�`��k♆O��<�$�Ov�l܏�z��8��kסf Rx��4�ҿ��G�U�_��w�p���桢f[3��^�����k� �ө̱�.,���Sö�#���ܙm����Vlp`��){t�M����U˷V�?���{jVsbچ�����9$��,�V�b:��� ���O�E�xнч�,����
:�S���չ@JH9�L���l]�����e�6��zv�|�O 0s]�М� <��Fܠ�BL��L
��X(l���Vw�h�H����$x���(4�!��y/XwJ&큋"PT>ɃC����sIF���A���4��5A��#H}��(&��
�B�m�<P��%��0^ؕZ��<��Qnt�~sO�K�+� \`���<s�1�@+��Z�s:G���D� ���6��-w(u��Q��֕�'��t��lJ���a3�=K�y^ �O�;r��Q���U=+�ٞ2�ux���p�]MUg�:������wo�Bu%�~�lû�LK�Z"EH��$��#�
r���+����S*!��,��n�{�o�
��P!ؒ%"����F����k�X�@�m�(����~�mQ�o�{�N�D��~�(��^�&��E#W����T%*��;4��vLѝ�Ǜ+�$^�ܒ�� ��X��Vf<�M(��\牡��'���=���.Ӣ(� �^� �!ڦ�Lo}��ר�l�О��4���ç|�(�A��`k�F����xX��[Km䁧Y�4\(��+��~F�	!K����/���K�<XTG�>����z�� ��<��&�[]�Ix�>@�z�Nzz^�'4*C�J��m�g3_Ӝ �/X0;0��`�"d	wM®��W�K�>�Vj�����*������b5�A��!�\�4<��,�he��袋��ME��o���̟܌/M�ĉ��bdHG�/@T<*�
�Y���ş��*�Y�MVcRzWTU͐�jbvU�]�ή*�xvA�;��1�|l6��g<��������ݺ� Ӿ
�'丁|0���� R)J���r��oۘ�U�Yqȑ�Ņ��� E������8Z�����#G���a��qq,
�؊�:VT�uL���<���(���r�G���x�"P�ci..њ���T�����F��h �#ѳ�"�����)h4�5��������QBr����l=�b�ZVhЀ~nqN��g��s�Y1��G����Ǟ��r��qz�S�E'Z�^C�!:��*�`����^]�.ws�-QT�z��8��r��G~;mFj��J���^y�(�ɑ&��&?)l��h�S	��;M�Ǜ �{E��Ɔ2�@��Gl��44k�1=�s�۠��%����"%�4�$j檙��SM�%@��ҭk��{����r#��Ԗ\/F�����(�퉔ܞH��*��(�`5��Kt�3	_���A�O���O���L�W���y�|GAm���Qyv=�a�JZK��,�ܨ�S\Fk�6�S�s�_PA�T��kUo[y�L�@�$E2L�	ț;iPM�Z(�!A���ДҐ�K���d��s޺%������U�OP�w|�P�ҩ�?X�w;�;���ج�ţ��t�hF:��%SR� �R䟸�H��]A@��d�sl#2ى����N"�̱��7�
-����'��%h��ˢ䱕2*�o׀����c��Z�2���.���E+UQ���R+�
[��PC{�b	�V宭�
xm�~�V<����j�Kd�pn��%~[�z���[�������l�L�H��]^6TV!�l(ݴ�(b�{�}�Rѣ��۲�6$��P���(�xd|E�V$mQ�V$mQіv�X�d�������C��!���x�p<d82���v<f83�U���?ׯ��*�Þ�J�Bb��6�������+��RX�*�ռ�ˏ"91��_��b�ղaDlR�I�p���)��z����?se