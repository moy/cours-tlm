XlxV37EB    50e6     de3x��ko�8�{~�..v�I%�vZ ����<����a!(6�U$C��dq?�f�I�,�vq=���r���������O����=������#�&2�E�%O���ڤmY��XGo���:�v��[2#7 ��s��6X�.�>�A�%/o�h��%t�,"��H4�z]�* �p�y���|�|/xn�A0> � '�O@L"��N��:,mCg�O��v$�����(�� 'O��e�L�4G�<I��s�>�Nc����a���w��o�{4*\�6�5J�3�'`R�,r�,��0Rb�N�#xqF/��5tC{�:ܷ���3/�)�-1x�>z�L:xB/�����'�%~����,p��C�^���`7����k5 ��_w[��M���_=�*U��$u����/
~Fy�*P�s^k`pR2�S/����i��o�\�j�q�&�<��J���:2�K�Ƌ(u��X����^��)y�_!(�5��7�>[_��g`�l;�b���+��"���t��z$��fQ�ާU��(��yH&�'�$��p��	��Q��y�ڄ>yc
��UP0G�\j-�b�Ccr��7/y w�9��nL5lQ8�qL�a6��W����T�<�`���r��^�n�8�����]�>l<T���}�F/dpzz��a��d����;�}����}m0X<��90���X.�q�����yz�X��r���짏�[�D�	�4��٣K��&�D���iJ�.�b�9d1`����z�:�cߍ��6��;�lʋwҰG;h =�&��No�s���������_]1�r{���,)����%�$IH�ޒn�lv��
��� ;`�фep�C��	�a�S7��Wg�5D��"���(q�ā5�a�ٰs5/%?s��QX��]�A�N�p^<�jn���y��5��I��ݔ��aqY <H�Bߊ�_��3�jB�g̘��޳���i0I���g9���;�z6�/�!�.�q?ѝ�[Z %J�Ȼ_�V}>;���F�C8�uT���۷�Sw�	�����D(E�yׂ׮�"��9)�! ��MF�ґv��av�q�`.���@" Q��;XLv!���:0k�+���/��o���>��ӵ���x�rЮ<��
�)F�5I&2�������Ke:�ʤ�+���F�\2v*�/f,���|5�})\���˛i�"Ɋ%�����S��	�^�)�����X����Ě��)���T�'v�P�|�t�wZ>�t�P?�9���T y���*�� ����c�*F���-�HYr�ղ��T}9e;{�&p"�?��ԄrS�ЯG��Uh��Y��ěNIM ��s�ċ{S�j��ư��T��b�o�+;87�)�%;�D�σι��24�n�8���O���&�
d+�>q�=��"��>�sQ��|F�Ai:��" ��^0s���WxS�H
�	�������A0��B"�!����`<���"h��iy!�ư	���[����J͗����R��waW��S?0&Ob�T�.�HI� l��!���3O���������LG�5�ϞO��d^�%����Y���ħ��LQ� ��(�"7-<���-�FK#�"#dS��%J����
|����K�����I��g ;��/\����Ϙse�������7Vz�3Q�a��@ۑǧ<b���������_cMŁ��d��꼩��(M�e�bq��K��a�Z
dkB[�m1?��I�N�K�DY|!C�u��p��F?y��Ά+C.��-o���=�e~f0�	�@��n�� k��5Ln(Bc��1�=.LM���sI\���C�T{�2�����hJ�T�j*�*�+�b�9U,��0�R����P�h���
T�N���=�}U�PAh�M��W�I���op6�[k��Z����\��!4 �TC�+j�/�q���hq����2i�t�B1:�ROr�*
/d����(�E,r����| �kj�Z��2I�M����
Jh�v0�`K��1]�Z�\Yg
tKS��,�\�ĝ����vv����#f��3r��8�~�J;4d0���?��S*�,ɚ�+�@�#�R^�COf����ϮJ葧�����
#��1��
�����[�f9?S��qH����[vH*�9������	ɜ���S�3<�P�=V'M� �Sd	vw��F�K����r{ҡG�'+��p}���I�gv٢P%�{�I�����5眯�;G���C0�h��l�*3�.�z�e�tZy��6�Ƥ�:���IZ�j�^�ziWF�o���ƥ+6�G#��	DW�~2��XIu
qs�w z7�$��IXf8!��6��1��凔T��O� ��:��*���n�ѝ��+���1H�U�T�۸��K�1PM@�D�Z�#����jS=��Rm6��qa��!~7��bՂ9���w�*������2�5����jh�Z�90�n5%�FK�z���t�yQ�QT�,~���2����Ws>�9�j����b���ױ1u��Ĳ2}2�v�XZ�xW�8L�!+�9h�ڶx��X�e��ϱc)hI����։W@��Ր�v��$E���%R�q�.��k��:l���U�.�]F7K�.��{��݈ܤDӒ��)���\�����f�Yx����j� kmS�b�j��S-�`�ƀ����Yϡ��$c{�{�N�JDI~ƥ2�;e�x�NK
BlGY8V��*f�����g���s�^��##���b0nf�k˔�L�u�qiI0^�D_Z�)������,sx�kL�߽�3�d��w���#�|:@6D���I�v�bؖe._m�䆥9��$���ƱT�['��p+�@>sޛ�Y�����:o����Vi��(�I{� ˍ�9�OM6�s���Vk��]ɡB"ԘK�t,9$�B������Y/�׽I�B���L�5�z��� ���b��~-�C2�[d�u{=~��|]	�wIW�$���Ky�3}���+�����b�K��%P��R�}�NuK����@��}�ITwT
��0��*�CY{��B���dy7A�+	��_��:	�_:	Xe�ov���I�uXr�0��Q������뭐�ˢ��m�2�n,���*?:�ꯗu��˸�+e[�5J��eY��2��3��_	�4�i�����0Z
��W��O�qRX����u-ǟaw����'zʪ�F��)�l�*A��>;�1��@E��lլ�Aw�����к���A��'�E�@�'���)���:F�9�^s<�W5G�9�0s<2��'�i��L����,`ݽ�r�1Z(�7�ڲПeH�X��[t"ڱ
�pۨ-h#����W�d'�ڥ9��.�ː`��r<5�֊�֤ز4�,�jc
0L�\ ���55�"�}�9uԖe*����/	�j�-o�%F���n�m9��͒�t���,��f�*�nb�&Ԋ��B.���&�