XlxV37EB    275b     9efxڵY{o���Oa1+�t)mg�^:3��ɪD�n{_�����	�����c;��@���є��w�}�'9:��o.�xh���e�h��C��n�^�ң���m�P�u����O۝��O�����(�I��k�~��vF}|-w���c�?��YL�x��D
��a�U@� \s6���y�m"�wZ���<$�4�|Eݖ\��-��C�Q�,h7�C�O��G,�3���m"�.h�p�ٲ�=� �F(�S4�����m�ǔ�ƨom=�>Nv�t����X<�>v�[��kšY��/V��(����%#�����D#\Cƣ8U��6xC̟�y����������E^��"6�uѶ�~��z�r��y�(��=כ�v��C���k]�JDL�f�)� ��^4~F}ʙSU�>>4`K�S��)��uH�O>y$�Θ��d�S���X=�n�YT�s���9�@�8'X<1��+1�U(J���YH=y����g����Y�� �����-��?>,�$�'��`�Qj�cB���LQ���e�� j��cZ�KW̡pH���S-��Mo�KF��h�G/,���0��!5����QD����o�����i��n ��	D'QZ�L��#�f�/������<U�<��	_#{0�� @�V��f�������<c�_.D�a R+�k����#Q�:��6&
���%��G�	'�R��lAЫ�Ø���LĽ�"�Pl�o���k{�s�����W�۽]T�dtT,�ey5j�Y���h���>��Mz����@�QAYr�4(E3�NQ�ϧ����%�Io|9����E�{��գ̅g����Ql���l���*T�@r=tT��W�����;���..ƕl��U�HK0��D��=�mAdg���e=�+OA�Q�+���8�q����|+�v�G�v�K?;�#84�|sU<�}��Bœ��=��-�� ���x�-,j���ci�r辷3�ǔ�kCl�X���r�s]^%�Đv;L�A.�N�����8�&�M���E�P;�K�����j�v�6�q��#QVs9�Vĺ6��*��N1c��A�hƨ��3���C���R��׫���? Dr5�|�F��oFY���4���EL!ԷR�(��R��>�|� �Is���EJc䍒�ɣT��%J�dd�2.f�(�l�Lp�0J�hd�R#l�Ha"ʋ�-��?�K=-����L+m)D���M0+q������m`�CS�q'w�'�I�(�@��i��T
������D����"
�z����7��R��w��y��$�s�~���QM����tЂj�֩�D����%�PdML�8���e
K��6D�Y*�aB��"� �����T֗����x��~C�$h���9���t�J��<'�`t�9P`�E�=��M� *���E�>�<]�D^�d���W4�\Y�����>"�D?��a1�rH��BC�CW8��o�B��l��m�Uє�.��M�\�4㡨� V�E�<r�{�Bxs{?�6�k�F�8�/�3}�{��(p���Ӡ�P}M��Y�V��T��wDW]�/���*����J�����$�� �����,�k�.�G"�;lӣ҇���\n^�T^z�5�{ڄ�U3��1�k���GqT��PX��2<pI�9_�:�NA�C��Ͽ7~���C"�:g39��&�3wJ0�M�0��3��͉7E�� _ءV�eĕ���F���o���V�y$w�����Q��y�M%�6�N:͓vF��rT�5
�����npds�*5�Ň����6y\��� �� y�2��V\y�
�CK���Z�R<�$������[���#2 ��1_���4�D�߶�ȇ�ÛHsܐ��4f�4��a[��-g�E3���=7�o#�п��_aN(����J�9� "�s����*����0�q���_;V�lW�t�V�<��&�v "n���2�@��D�&�� ��I�A���Y�+sP�q�,A�s�r����2�&<�1�(q��p֙�z�4�$�'m�Ǻ�{c��X��3���M,6������cJE_`�J۫��o�m�n��7�m��5?�T�7#�a�����g|~?���H�Rd���O�H�?|H�ϥ{¦6e�OT8��׵t@�v����7�p�x�1��4�L���uS�E+}+�9��A\Vp�Mk(�=ز���0�4�pCgK?yW �g�_Q� K�V��E�r�i��q�#�T%�|Ë/�Cs֕UK�
�dH�UʄVʾ�!�}g�_�i�q#�|=g��Q^���7���Q=��s��Q{�l�l�q&��䓦;�VH�nY
�ԲSU��M�� �L��4�è�7���F�,�]V
 '|��z5�Xm�R�Z�o+4)���T}����>3ֳ&��� ���9�V^�v��i\9���S��8d��X�V���N���M�2-���çW{6���[�Φ�-�����﫯3�/ ����)