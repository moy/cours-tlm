XlxV37EB    7307    1225x��]�O����_1J�n�*P��%K%�I�R�ޫ��I&`��Y���?��Ïyڎ�j7Jb���9gΜ����޾�}::�1�gr�ik{���5���֛'��xӝ��Y����-��[�~- ����o��0r0|\�=7���S��(H���Mo�M�e���Sү�yS�1��p�y7�	��|/x�q0�f�#�� �Qt�f;�N��c8F���d<H�B�������	��;��[Q<��E���-|t��$�̗��܋A����<�XL+�f��V��^'ђ�h>���.�9��U%=G��6�
���I�|��$��clƒ���޶���yQ�dC�y:���Ҭ|��;/���*�'��>ȕ��!�G�@��� ݧ��	Z9���?�	������?�̻�}��*ƛ�٤��0/�
P�M�H���#[bOfh�x�$Od�|��|�QƉ� p���t�	�t��Yl��.��La��My�ixw�.6F�T��]x�.��|�#D�4��w�L8{%t�H˪1i����,����Q1aq�y�7���"\&�ea��t^���{S��ʇS�6�Z0f����9(�Xsx�[�m�@�ԍ��SǨ
�q~��dxy)�"�����	*�2<��'ߝc�W����|ظ����ȍ��x8����v�d�ܰ�n���A���7��k��9�}ǲ�Q��w�czi|y�p��N��L;}�xNl����Y�۰ZYP��2�K8[�9��[���-2�'ηˡs~����]N.��C�P"|�h�R}<�9���ӻ ;�e��B7@��`�O�zvF39��4���]pFG_Ƨߩۣ-���{s�G��9Q�;�|��}s.9��	rT�[4�Skj�`�^��S�t�uH<q�g�,�G�0j[D\N)۰3H!�u!�8��Q��D��}]W�x��nU+�,�=�{]g�� �󕴢"|ž��2ə�Lƌ�$���1mZ��)�qq�⥟�q�Xy�f�
�.�	o��0����jG\V	bD�������e��������}�2���`���x�G�2�>^��^�\��L9'�sn������t���Ε�N��2g���T����S24�"�Ye3��V�ɓ��LV=��q2kf�8��Y�h,5�ܑYf4l���L�E�/I��҆�����ح3�#�W4�1�]�q#�!��K�y;C�E���a8v�Ƹr#70y��6+?�
��͜Un<E_��3�yA�Lh�R����B�0@4(w�5ТP��Ti�0c�ش`��zև��|3�����t
]�t��n�H�6��ĭ��Q���0��6�q<o����f3��HŽ���t����	w�9�1��u��-Z�f�.��/��5|nQ ���A���:5����>q���'�Č� �\�k����T ]�$L�z��(b��tZ��vq�K�sWJ�;,����&�P����.p�0$�)�eY-�����x8pw�M�h�/A��őHE��Ե\�4P����AhNy��MK4�u�X������ǐs$�L��btb���+3��dP�H��솺Of��zIF[wgK(p��n0����*���ii���ލ<Ϯ��c��
��Ӑ�Cܺ��!�f���X�*O^嵋�£�H#{�?�O18wc&�7m~1���������.�I#b��1@���i���
�a��9~֜ؖ7LIL�a8L�ƕ�pH#a��ˁ{�IE���}Z
�j {�%L.�(`E�1_+��g� L�ee�	���ь�YQ5ݳSM��/��1�rK�ҬT;�kK����)+D,HG��TV\���*�nO���_����;e{}^f8	&I4��}?| 	� �-#��ξ�)�!����[L�����1�"$��;�6�IO���� �=� �~vvv����}�m� ���h���k��بgu6>TM����)`��I+÷��br�a�#]��.<I�J2�16ar��|��["���J%�cT߽F�z�
Jf�,#T��J�������sy�)��x�e߻�����I�LRk�{����!�9��W*�U}괒�����6-�ei���ԍ`X��6���& �*�������|I�� H�;�zO*����Kݺ"� r�Q%��8DE(.u+9�,�R��RV���*F�C��U�*-�B.�i�L�,��
20/Y(7�7�* ;���������9��i|�m9*)2�ڮhy,_�
Ơ�+?P����cF�5��U��Yi�,rή�=�j��ݼk���X�U�������Ԟ���@c��`i$YS���&X�u�"S�ʲ,�GBȊ�+,8}�Ɂ��9v[YH��9�6��ꛘ����hJ}�_�~�*��ϩ3�0Y���$]q�l!��(�s-��4r��;��d���ݝ�lK�K�1`y��$�Wj�:�Z�#��
�UGR�By%U�k������w�9V�ݢ��,I�I�8�Ⓡ0?��|%��R"f��z�~{�^����dx��ȹc��8��Ь���F#X��5ǲJWS쎎6�y\�Z�\���豢53�dy#�N�^�F��FAݹ�)(�j��"mȎ"�er����d����P��a�?�����T{�F7(1U
���2�f����ݎ	�JE��#���k�E��_[��r�l�%䲭u���r�/"���\v�\�����\�
�^�o�k���eA�n�s���-�AE�8�c��d������#"�Vs���Ҿ�z�ݪ�64�ݯ�6l�6����e�6��[�m�1�b߭�Ȫ�6\�H`c#����g��^�H`c#����[��u�66]߭��ېڗ�i���~e�5��3�d6dX�7��掲��֚�s�YIM�Jyjⴆ�d3N\��D6�!��&d�7+��!���`���0�5Sz�*t����t�Oq�G�T���Ȓd��J�҅����x<�C _�>~=�4w��?�[�O:�Bw��.��y���m�]�,��V��2�)�^]q��e��nGv�����l��gN+�A㎟��gt�`�m�����ӥ<[���w`åV�7�
4��;Ȋ)�u��#=)wµ�ϴn�N�SL����tj0w�g5��f����>=����}-�M����n72���j�=���+t?����ov���~-�M|�%�����?���74������>��ܐ���I�ￄ��+>��Xg+Ϊ�����G�n>��>9��gJ8h�$l�Y�r�O����,+���$���B@�ѫa�_Z
�,��V:Q˟��Ԝ�e�*��I_��	Iml=Wl9��Su�����ܷ-�8����⭴����n�F{!ϩѾ�+������4U-�'��^Y�t[��j�j�e0����s�����%(�}�z�j�
M�i�����Ҏ�Pk�_�FJdn�j��� ���h��J�������$ծ`�bC������������H�R[Q���5�'�=S�0(����E���Yl�ϒ=� �tZE���Q$܈"�ϢH��"�(�ވ"�P��<B�ZA7[�NW����0B����H�障'��H�J7D+����z��j��\SQr���@a�[繵�v�V��׾3r���c ܬ)¿������uF[i��L=�Ԋ�$9��������B��X)���n�Y���E7�W.��뢴�ݧo3��;���:����R�w������]n�no5��
������S��S+8^	�}��W��Y:{5����?���^�!�J�՜!�r��%�C�V�C����ُ6w��H�\F1P%'���������V-nR`�ĥ������Uϫu�%gkJ��߳�W�-~��srbr�(o2�j�WS���1����j���DS��Q����y�tj���S��[�,��org��!TO{���2}v�)���{
}~x$(~���
}�����#��[����{u�ns������C2?��_m��W�X��e���T��J�,]�h�Z{g��ڣ�`Ru��"���v��%�c�]��)�6�ǣ��]gK�0E�DC���["�$M��+�G�i�z$���� �=�m(ɔ�#d��G�y�vD�����z�2C�jB�pѯ-�Dn���3�i�`6pSe�.��Qp���w>�x����y�����K���a����V�r�16t���a�k��tE���o��w7B�KL�a(�漫����2
 $(��,�T�73Y�{�
�`5`���ֲ���?A}�7j�)	����
?^:��U�dH�oH<c�%���!
L�!�{0E6���|r�H�����Y�8��Q���'[�H���P��P���i�&�n%�^M��J���H��H�6oWC��:��%�:������*��'ܰ���U���,�	=��y
9�T(J5�6�2jey��eAy�����ڠgy�u=ѷ�{1p�KxI9�<&�#.6������9½U��:�*��w#��������m�