XlxV37EB    343d     aebx��Zms�H�ί�r�.�؎��|�$U6/>]� ޲�jK5�T%	b���oϋ�i$��N�6h����������غ���&W���� ?��5k�uH�$v��t3���t��o�yj��a�0��&2���[�'�8�p�����B݄���d�D�؍wp�,ݘ8�&$�01���yW�)�N�ޅ�b�;�s��cd��)*\xb��$"��N��sDz�%���4>C�~'a�~J���a`:�%���8�Vk��`iQ�$`�(7N�#�\k���r�$ �j�	��*���x���"�OG��Fq�Z\8��(5O���#��a'�J^��/���-���Z��0�� /��"w�c/j!�����(���j G9���1�g������ǣl�hŇ0KQ�d����u��߱�I�D.�����wkR�����'!!���0�7� �<��QKc���l�S
8G�9�j��\��^��(.XI���&�/��pG���w
 ��(n|J�oM��9~�.��z��SA�4�Kgb��q��9
6�z�u {��s��fd�:����P@#�x�����!���|�Í��v�&��#"q�D��ĸ;��X]�u�S7 -bщy����{�kro���o�ۿ��|}�TQ��i���z�^�¾�F������ئ���{�4�oV4�l �#)�o�S����s�0l�a����%{4��(8���!^�0zd;�ƞ������+Ζ�H=Я�J�C=tF�|�^~]xAU��ܨ�f?T�Q?�@�9��M�i!���_|��,��y��9�[{�c�`�ݤ-H�b� aBs���l�8��\ڗ�c�w���L��u�g$�6��N��=(S��+|�O8b{�L0�`�[#�g�
��o�@rm��mVkT1���.�qoo�dº�� ���u�78�߱��l��2�FLFå��܏��
Z�0r����RLr1���\b-��ϐ��ۯ�R��"��ڗ�b�Bַ��iB�V�0�c���
�i�hӺ�:����ll��n'�<M�
T�b���	0���X�jl0�'A:D:'K��8Hͪ�f��Y~0������V���=�K5<�j��U4��Q�YT���`b_\w%E�=߾�a^)�h�L<��]��pє=����������Q�H��y)�8�L EP���2BGPo96���:�Z��P��B%ؔ*���槞V�N���]T:D�����ua�5ˇ�J���Clɵ�0&'8ؚ�R��'��t%K'���5�fCb�WV໾.��/�~y���j���0�;�~Q;��è��=v(ퟐh��Y����f%:�\]g򺮭�up-\�\��#"[�$%�d����6���S��DV����YmL��󁅴*y��Ff	=�k!t8�e������B�	������'ZpY[�y�h0��`6�G��i�N
^��.v�.��J���x�eEw��q��.�p������'8\@_��k�Hk���hi�0ep_O1��v��b߆�g�6wE6wUl7�i�����U�� T�lT�|�$����g�g����'�[�r+�y�8�x��}o!��E��1�A�,@~#��s� ����M;����	����0Q]J&L�DrcM��d��U��mb�o�.hʟ��3Ї/h44���c¶MV)$8Mf֧t��Uc؟\+z�Ȣ�U�1���6�ƶ��G%	 �Q�������{�&y�$<�F�yb5���I ����eK�d#�锬Y�uZ�$�1L��p�}����J�].fvpU�*�iM�=�����z�{�g�zSC߬�oj��
�3F���l�a�N�EUJ�?kA������4j���F*ma�CY�!���+�LmI&�%f���Z�;>q����X�eB$�3S�AbdyX�9+���\N�a��W��%Y��' y��#?(h9��RM�ӉV���Z:�Y� ����O(*��a�&��Vʝ�I���P�N��<{ׅ�G�
;���VrS����2�Ǻl)�|J���y�aqh�g٭;.�D�����%��,(�_��V�_�[����e�;�mŜB�|���n�Z���J�cK�wg�l٤b���> �7�d�R���A�*�M�x���ߴ����R ��r���7��V�y��=dM�f�J����)�Z�E�<@3�d�~w$\iT+u��"�p����J��@���zC�UBG�nT�H��/e�R���04_/��rAo��t;Oc�6{�N��&x��l̏��>畩h�n:�k��4M��͞��fo��pP�f�/;[������Hʊ�4 ����� �-���X���խ1�[�Х+��L�-H�uty�{~ސ3��Y��͂>]S��Z��t�D� �>1ӊ#�|�f�Y5��i���)ڝ'��_�{��DRM_�+�Ł-.Q�7>]]2SSg�e�C:�����K��7�$WJ:��F�gix��܃*S�.~�ݩ��c;���%�R��-�	$5�P\�Cu:�8ƞר�v��"G�a�G�x����W�L��DAbOh@��ҳ�
q�f���a�Gփ�U�8��en��ַ���)��	K"�G�P+�:Yj(�N�9܋�ˢ�����w�a��H\𭋫�Kw�lHu�la�H�;}�g� s���ܙ3�� U�����Зy/[.*��)>#�~q�Q~�J@�!*��LO��@�К�J�vy���m�W��/���