XlxV37EB    3f74     a5fx��Zmo�H�ίh1+d�qBLF��Eb�(�=���2�CZcld&Y폿�n۴�m3Y��!�TUw=���E�Ճ>�j�֛��|��j���yZY!\�HU��'�?�*R���i[i"��]Ww<�}Y��
���jh�2�)�\b�*"�G��O�c<S���!h�S����7���'E ]ًW�Ξ=4�&�^*�g5�.pa����!.qVdZ�}T:Ʊ�P�X���������c��8.����pMQtF�&��Ѕ��u��C�$��$lY�z�hB-�yEb�)�=���q��YrWk�6w����C����l;kk��Z����%��;u=�ym/�CYG�`\UU\xn��z��d�V��t1e�o�1�z$p���Z3�k��ܶ�vhm��� ���\:�t�m���x�Y�P�0m�{���2���
Ѧt�!x�᥸>p�^����lx]��3b�kY�B�J;�Ė�Д<Q�{]�t���}W����A�+-�,�≯�	6sS匥��q$���!���*� ��C19{.	.肘�퀙g�����F���ȆK�qn;��ay'q��ƒL�0S�H�Q�0���d?!{�-�Z�P%9��mJVԀ2E��)���kn�xx�M�r�H���q�%�j�m�%�V5��A�h��� Px:D�.4.��{;��ڗ����_7��W_�*��{L:qX�ѭ)�8��s �^�`�^����n�]����iϨ�a�l�t�섬�u�\0��Q�7j8����$ڪ�)�����k��K�Րe�P����Vj��s����5K�����k��#��J^<|�uh��C��̠:<A	3_+�$3�&ts	q�;$�k��?z��{�x�롒e{HOt�*�cz����Ơ�+PO�=�<JY.  ��PI�U�֔,���m
��LY2�Px�t</��qL�Q\�Q�"��϶=S��~�$b~��bp������Ԁ|;�> F�	z��]���ofY^6m�k<;���?c��A����Ц���	�����X��*`��e7&3|x�_����V�\���>�<����͈���(����Ʉ�b%�t�(�^�xQ+�V�E}y�����eJe�+��D�@As�}}������r���1:犔Q%��,�	y��i�/��Ì Tr�܆�Y��%B�s�k8�n!lQ��Dm$�h7�z�1�;�H�h��en�>GJ@e}7o�هъ�KN1`�ݫ�&�m�b���8�̸xo$�=�m�[͠���m��@� |Z�r�+>�x���}V.)���?�[���|�(rFǨ���8u�����ݳH��ΰE��NW�iu�<~~��`��y�I�%ԓ����{p��ۯ���0��ú�<tz�<�n{��'�󏈭?**J�g�=A�8��Ϸ,����I��5N�{2��BHCf��S��M��].X�k�o���Sa��B�A�K��D�A�h!��sE�s=��h��c�!��u*�fcb�L�Y��ॡK���'���}��g��9�8���\kn�3y�J��D:�ig1H����p�	�%������m���0F�6�/���[��D!>GX�O���f�����vć~���F���"`#��ʋ��Ő?4Ct�͚�6�~����s���T����}A?�(s�W^?��\z����?�~��z h�p�b%�+�4F�ش,h�<Cq�?�vݕ��Bp�>�J�,��]��%F`�{'��{x!� {�E�F�̜�t]��
����+�;QN�3J���Br�'{�	�)s}!ۘ�2��.�����=OZ �d1��@�����ٿ _�[^\a\0�ɸ�a�NcR%&L!3��D833��,:�ӛ�-�q#�TX1�Ն^�h���+VDƍD�滴�I»	���ө�oeiB8E���+�-ͫ�v.�ĕ��̌�˨()'�"��v[B�
Y��;�,���9�����)�wJ0o ��?������RXIȫ1"��!MJ��7i<M 1��� �&y%��/{���wq��d�K�2�X�������zTҸސÒ\=An܇�'�C*֍Zb�����%��z�uIq�`U�S
8Ĵ�Y�RֻD�9���L�G�R�"��~EV�"u,�m��E񛖰׈0b�g0�2�h^6�1�K�s���k�f?��ś���~Tl�H�R��)��L��8��ɛ�DF?B����Մ�^���-�'mm����ܓ
!u��6!)FPe�X��+��`%����T��T��TŹTm�i3���\z6��W���S=�{�rU=������m^%p�ց���yW?��{.~	{G�mc���,aw)u/���RIY;ar�&���l�h�gZ���%hsb�������Hs�2pQb%y��f.J|��.S�±�p�^8�N����^�&�o.�L����\�%�#��&+�D�,UN�]5R�ꙓ��������Us�Y]c��*��g[f|i>�2b���okT�������lYy{�2e�Y����?��T��%&�q��?,�d,G�_�5Ǎs�����ռǭf���#����ڣ���L�������1!��q8,� 8�o� ���B@*�~�*06�4o��7�Û��p_����-6������N��_�<�