XlxV37EB    80f5    149dx��]{o۸��ߟ��\L�"I%;��t��vZy���6ًYA��D�#��6��~�=��(>%ٱw{��$Ϗ�!y^<�wv&�ӏ�#�h�M>�v�� ��x�'��Y�����E�yw~4_�Ow��'��8{o\�M�K�n��۾󖤙��~�����M4��4��􉶉� ���������,�e�I��ʱ~�y]�Xȇ��9	o�2r.���6G�]b'8X,%HI�A��w�U���a9
A�������e�#H�0�xQ���:����A:K��f#��o	�+���O��$��0�%������i���%���$K�T�
���D[��8)YJn�ď�ͧ0����H?&�v���K��0I�bXX���)�a��v�w��I<o�`NN���cJ��^�$��u@��hvG�ff��hEq2�s3�xrH��#�c���'�j����A���>~
�a<9 �6� 0� ����K�"�}����eáV�$�@FeA4��0y<ڤ	�%��q��;�ϓW��&j�m0���]�����ZUgE�m�ꎩ��ᔽ]r���Bn�D���@ݜtoWd3c1Ԣ@!����u~�ޅ��Tl�i`���r9�����φ����R�C=�>����[�ϲ����A{o#�����z�E[�j��g_�	�l�uk������/��|�*]M�`1" ������A�mVE��?x�2�U	�7a�����{>��<(A��̽�A�F�����o�Yj��=&	���f"�,��#�U�/*�t�@�>�?��Ip��y�?K0@8�E��1uc��ze��i�d{164��6(L�����?f�y��h�²�y���dT=�@eD� f�l���б����|�;r��$3�H��ĳ M�:Dh�����Dڇ8�i��ˇ����>:���W�c��_�>�8����EEk^'~�Lƣ�h�B탿���[ķ��s�w{� �/}0E��[�tΒ�z��xO{��x>#�?ߥҏ��0�!�o�}�Z�^�-���Ɔ"W�ixϪd�W�F�MH��8���l�'ll�?n��7� a�jqI�-�L�9:�8�J3�O؇�������ʼ-n�u�M(�J3j�*O�=�2�[�jxu
��/&�d�����u/�{T(�2��F�w��Pm ��[q�3�f1#B��x8�$��$~L@X�1v���w{H���L���t����T��ô�J�f��W��9ՠzɜu���G�8��;�J���b8�H]��\�.t��z`����=��'m9�v
��
T��kD%������:]��L���ɀ���hÉ2@di��C�{Ae͈i��6��F���Q
;�;{��Q����	H�9�K��F��D�e�1�pͲ\Ր��g��l��*��O~"����u��C�x;���P����8��N��H�t�)r�(+BƧ�)��0�� ��!�Ԇ{���`�:�fd{3�Ҝkohcq�\XC�������*[�����R8
N_��/x��_���BW��*�\Z�亸п��QN���|�����з�oR]�����o^���q���1N�� ���5�F��)���7@=�� ���\mp����k68B(�\�p��Y덣:e.�7N5c�0WoUpuV(���b��p�]���1/�x�L}?���c�c���k}�k ��Cb_7�P��2G�[
�����2��W͎�2��.Ɏ�s���nu���}�:�$�I�-f�zc*�K�3h�X���*�.���"�Zj����	��H-p�hK�@�l������o a-7a�_b��j�*�S�;&���:�k�V�5Vb�pU3-�d��ea�Q��_�4�{�2��'��5bE�\�Lˊ�M�����h�T��42���#��ɫ�'��.��`���#�GH�a�=��[`��?�����l�K���#Uu�z�k������jt���߬���w0�{gS�xt4e��Z�NQ�>�������O�ƵT��4�װ�|���@��Plp���{��}E����4 ��W������[D܎��y����F;� �s��v�ҎR���Z��m��'+�s�h�g)(�����Tn0r��oޓ��q��N~���I����s�$e��=q�)4E%4.�)h�J���h����Qu����XsTym�;�ri�Ԡ����@��Ч��0���w�?0�V����۽���P�ڥP�ۦ�B��s`[�����JD`��%�`���B�ih��h�HC۶y��@ӣ4fk�H��\�5���]�����e��B� ��0��J��,GǴ֋�ͱM�<����{Q����͈���˷�sKY�(ZյE�&��_�X+���ZB�6�lDZ�TU?����\iDu�
ꊤ�%&M��j�U-���ن���b��K����	iC`�m�f!>l6�I���Il�{L�a��-��Dh.��� �1�4gFnn1S%M��d��7�x�qv$)
m08;B����pѿ�)S{0K���f.-	Ir�D���u��Ӄ����tr�|��m �.�m �]�� ����;��b1x���0&����i�~��Y"/���y��Ц�OKX|�{���.�b���Iӡ̖�n��ns�O �s�*�}������R`��̢����f��V"`��,��p��>9��dv���E���:��^�㴼۴�Ӵ�����ۘ�������f�rk��V�m���m�U%�Ҙ���8W{M���Os��i�ڪ��B��<�8EG���s׏i�����	��;���ȿ���Bx���m�ye\��1Š ��Ѐ@g�4i-��4T�(Xd�M����t�ސ1Ik{�v�;8磃!��ǅ��fQ��V�ِ�s�j��?R&�:��RǼ�����Q����WË/�c�'��pn�m�{~�0��NV���&�
�1`H{A�RS���BD���p���Y"�!!��V�!d�E*��U��9[ҧ��d�HS��<GFf/o�v�5V�0W:F�¹�Tc�*��C{g�pm�F�,�c ��e�z��ԫlK(�*�	�\��況s .��R�� z��̲���ƿ���x���`Q�$�X��ԇD7�bò7�=mѷ�h���f�k���Ɠ�Ҹ��cuX��AAJ(���`�q�_i�S*�h�L��eMQc4��D�cL63��y��t��9Z�N�$�f>��Q�N����	�u���"؁Cȁ[z�Nΰ��q�p뿏�����{n��2��K6��KnD8����".�'"9
�+)��[���Є#9�[��T�DG5��qB��m��OWݻfmʻ)��ѐ����O�䚷Es�k�E��\M�H.�
�]�;Udɴ��Ji��b�T����#8�1�2_�di�8�� Y�Z±1��W��DLVO�X���ʖ ���>����!�]n7���?���]�ބ3<�}�'� ���[��w�ո��R�x*�7�9|�_\�e�n��,g�s�F���h����7�t;��<��1����@�sVm_�$���<�Ah����9�.4u��k����fQ�HB��+�fK��K?���	� ��QA�Y�?�sqv�x��&U+�[W8/�7)i����N�c(���`⟭b��.�,#�j���K�[�����L)H_�8�%ʨ��-�)cg��4z�zxӞw�>�u*m��
�_
�}����x�����i��׍��E ���%ג�D(���U9(WJ���.M�����T����P>_a�P���P"�0�]��&zf�򭅠������f-���93�"$��]�T�24�H� ��I�1R
Xc)~B����-��c�<�K��~���/�^��ɱ�{3�p�fڜF�#�� �>ߚ!-N��d����v�鮿���[���(, �,t��׏_��E	��@��N��!S�l'%�4�"�Yn�榹�0�m�X�,��XL�t�1i��;xD���u��,@#Z)o'6�\�V����P�o�UGacpugG���#.h� y[������>ٔ��]9z'@>y��*%��]���]�����؃挫%�������s1��o��,GU����	�,��|>1���Ɂs����bo��#��κ�쬋�@�mt��Tz��я�v�,�§��X��D�^�o4/���]�+��W$�v�����xlC,VP�'���������e{��X��5�5Dw�k���ot���^�ɽ�)���������Y�������:�ނ�+�tݗ*]��B��X�j]f�Z7G��rk]>�)I%V,�^��%j�.�tMm�7)l@��)l<��.�t=�g=Q��[�������(�Ň��1�K�_�g(��@�ׂ�$nW^�Z���
ϱ��F
�e����*�����M����Zg��W��<�b^|��HF�e�Z��f$紖�j��L"�7a�7q�@v��vA�T#HH�-��!z��a�n��v~�r~S�8*^1�CHB�1NAlU��a�ngC�[u�D;%'�VR�,���j朥3����9%qN�����	��K��~��E��^�xY�8\ݑ��--Cʍ�Z)��r8�%��g�̫�:"˟Ϫa��v��C�py^n5hٿ5�������o�Z�Q���*���c ���\��߈���f
�i�ޣkq#u�@i6՗�4�:-Y���n|�Z�rɫ����U�f�pK�F�X���dyѕ8nx�+q�f�zO��d�D5�A����5R�v
�\G���\G�Ja;Z���Xq5W��5�.D)��a��z�e�R[��a��ko�Yئ�:Z���7���~ FhZ�����_���o>A��'!eNyZ���t١�N�w�m�_J��*�IsJ '��#�����/�.�C$gX~8����`�!P�BS���I*1&e��E�j�ե�Z�mS��BM72��T�sS$!^�@��"M�G�elN°(#����u¿йq�YL�H�dkq�u�b*O9ϏX��A>�cӢ ls˾[�bn�/�a�$����ä��<�ǒas)��'��ת��iʹ��*b��_sȮS�/��$D���>��m�&���L-��xv3��w���u0F���U)ﭜ�l�Ee���#/��;���A� \��t