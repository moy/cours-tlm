XlxV37EB    1cc4     739xڽY[o�H~�W�H!Q�@ڮ
m�lBT�n���}�{�Q͌wfL��?~��`���M�|9��w�$���^�z��A���#+��4c�6��$8�A�тv���e���݆f���u���e�0m���Q����u�I+���i",�m�y%�ӧ�Ry �*�k1����	���s�&B!Ϡ/�\�!8
��g<h�ꕓ�$WN��D��т��eB�����������c�X��<!GJO��h��3@]fD�aly@��%/��
�K�a��tE�K��a�!6<8�!�W�@���Ri2������X��IV��p�������G3�`a$kΧ2�)�d5;�}��>ȩ
Ĉ|6*�>��1��F_9~Aw���7
�V���2y�X�.��4�_&"!����g����s��>���<�UL�6b)ΰ��2S�z��T��|C1N�O:3"�E):_�`�(R�6~g>R+>*��Ⱦ|z��`&�����~����YL�X}|���I���@5�����q����p)d6���B'�猺熣>c��}S, V,5�n'�A���CD���D�qtIDNϋ<� �E�@a ��0a3N�M!���*× i#tG���3IR�4?ʲ�/o�����W���]���C^&�A��&͡�a���<d��瑟MɬG0���0��@tQsW<&��2|���XEMeŔ�Ư�����s�>�"�My'��dJ7�+n|-���ù�~��/X}�A��DK/�ߞ?��c��u�,��ѓ�rۉҝ���¡I_��L�E��:Z����������(yS��I��N)=�$�;}���v�uNR�����4�3y~æ4�/�����8�Y��
����`���t
��z���7-��v���ध/������hU���H� �A[��c.��6ք��;ͱ኉[#9��{~�����ġi�;�%��{�)��)��c�i��dE>?���G)�m��">5�1F"��������d^�(�%Q��I�ԗ�t�,�hdma&CyN� m�+���Ql����Xj�Iq�Dx�ٚz�B�|XP��j��u.C��L�Շ(���E)'M+Z'�.�h������`���HI*�1�fI��3������{�޻�^?�\~xr��P�I�[��pwc/Tc�{�֛W��J�'��ǽ��hJ�U��Kop���^z��wq*����{a�pGwҭ$�������К˺���I)u���J�^op��'�g�޴��h��I82da��]?������K1���?�?c�.����0j1���Z�G}}��AXN=�����~���T�"Y�����r�OL�e{3<�(]kҊ��$u��E�[��[)7V~���\�]T{)7��N��a��=kI��{y�#����n	�K�e&�!��U:���$h���b�C�]]_w2؅b�I�9K��cJ�#��cN;�;������1�>�[nJ��	*9�\��9Q3��D+�b��3�t����T2R���PSt�4��7��<�B��`���!ωS\Y���렺A����F�;nX�\x�
���m���E�t׎#+�1ʋ$�kD+�V��O�{�[+�.�ٲ8Q[�zT:4\���"zط�"�*ǥ��%yhY~�,Y���u���Б>�̢)G.�R�j�,����9U������ۜ���5�?R���m�h�o�rm��#�����Ϲ	�]Ç�zÝj��l��kݸN��ݬvK� �s���o5wj(*̃�h�v:��)��N���A·��`(]��A��|�t4ǻ�� �#�