XlxV37EB    15ef     685xڽXmo9�ί%���mOW�V�(U��4*I��T�̮�����%�t?�f��e���N����x��i��4�m8���֫��8T��\ĭ%�:=�w�Ϟ�zO�}��ϟ���Xf�F��4ڇ�h��@F�
�T������7�b8;�S�U��b����I$<��
��D���eԁ7In���Kw`����]-��o-DJZ&��L�Ln�^�ht&b�ı�!xBΔN�J��mZ��+�j1�-�����rs���4fZ��-�̔�`�!7<n݃�L��(�DiR&J����
�\��IV�]p�E��n<����%"��ds�y������M
��������Ōl6*�GbN���L��g��,a8Gdj��i�Û�2r�uKs��`2aQ�t,�d/f����]��l��E.b:0��Cq���3ma�Z�R���c��y~ҩ�Q��B���Q��Y����JZ�W�+H��{Ɨ`�K!�$�ѝ�Yt�}|ɓ=�>KnD	��K�ٙ���ܸ��Iu)a��	1Z��Q�\p���xK�MQHC�C@�v��,�p����B!�Ҹu��f�q�/I��(ɋ!��[r
o�)(����>���gdF�$�0in������]x��޿�йKݵ{��i��Ṓ�S���������u~�y���c��$+,�9*�&jN��s|_}������ʊ��������c�;�D�%K���<�5@E��H��B�/s�m?4�C�=)�����鋧������5c�]�l��x�ۅ҃��s��#�|�Ka*��9Y�Pk{�X��U>�#��ޓ��1Ք^��n?p��v�By'4F����d�K��*��>+Ҡr ���_�n��9Vf3ؙ!Gg�<�����~�-ॢ�����by\���c��b�0d� �uY�Ϲ�ZDw�z�axV�f�C>s%Ʈ2���o���$����eI��vpf��E���C�,�rQ].R�M%���Er*�	f"㉳[a�������:
���V�瓣�Hڳ��E��¤(��'h7�
j�6�Yn�59��-�$��"�+͝�G)\S�1�|\�`�0E�oL����[��V�8��Q��ϟ���dӵ��hb����~9��_}_�×������>x�H�T�ƣ�輁���:��a��"
{�ߟu��=o4��i���ֲQe#�{"��0 �\��y������>Ƣ8������X�_xDo[��[J��.u;�E���"���,����6��[��<��d��h�U.�H=[�����j
���E���%��6s���0<q&��=H��z�'�&F����t��D�چb�ۿ!�s�M��.����Hw�I6|6f�6-�3�A�"� �Ъ������*W��w�m��W(���z���"h�F|��~g�� 0�t������Z;�8G�����N�L�/
��iJ0����"�8��u�nd儙���GM�˓`�P��g{�G��-�<�l��Q�b�l�� �8D��_���ᘢ���XW]�̊ܧ�� ��� ��ύ,�	����
`� /)�z@o0�d��A0�;qd�k��jJ;06
���.���+u:���R�����o��I�s���瀾