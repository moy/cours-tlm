XlxV37EB    fa00    235dx��=is�ȶ��E�g�� 	;�$S��$�xI'N�W*��
H�$�L����nI�RkD��\3�Hg�>k/����Z?[;;����L����~}7i��u����ޛ��F׈ft��C��ܒ��9�uk���$m� ud���,�� �#o��;�w!��L��E��5�G�O��"ķۿ�'��U��	�p��k�샨�"��ƾ3�e@ʦ�ů��Ow���N,��x�ž��vC1>mx�E�N�ξ��<� �x����w.�{'�e�_�+�[�R�Z�} 6�WvE�x�r=|r���Xg)?��N{oG{�T>8~�����6��sk渷�	��Q���q���d�=���u�ip@T�헦�c����G1�Ol��/s�������vb�eab )$ ��-	���ھ3.Be�G�Km�M&����>����_}�|"`!h���^���c�.(d����P��X�{���Z`J�5-�y3q���)�烘o�i��֓D'�H.B��d���_����hj!cCm���� ��3? ���|���"��p����m�[�z�Q,@��Z�C=��$�'�#_�s�[�-P�vEh��ˋ���PV��s���C�b�F~wr~5��n�60������V{�ؚ:#��c�vo���:'�ԻuƦ��u^[өp�]���L bwb*g���FS�Oۼ��i1������!�t���)���u;��#�ݦNM��&f�p!L�Y����X��������H��ub�a���X��0��O���%q��8 ���ʑyl^|>��:�-8t�s�h���l<�f^��>�x�>����c����9��dYī��Ǔ+�����68�Nv�����<�O��Ǘ ���=���h��#��D&߶������i��S5
���)�OO/�#:חe�m�x�:��<\����.�:a�-����z'��/������-�U#�_̡�1*D�%j��l<�]@ܥ��Ȁf�F{;�FI�d��?�A'�c-���zg�yS�r!�pB���.���,�?��)W!9f!����d\���0�k�F/av�;0p��̈9 �mM$�U+!�-͡=�A�H�)� 0��Fvqgi?S�J��'�;a�JRifZb�{���BK"�ܖ�[������E`�ѝ<�0���(m|p�Lt+[t��Q�Xoi����Cbzf��H)�2N	�33�� Dr O$���7���&.ϯ�� u�ۿl����}��?�3�� ��C���y�3��srolڈ<�!��X�0���?\�ajOn�	��;�jW���l^��l���m�
�p1�2v]]�s}l�|4Dr���o�m�O��:vi���["�''���C��#L@���biT�(Ͱp���,7�Y	4��@1FTOr����J�U��i؋/W�;��Qʫ�t�JzK�)�k9���T!�hC�	��罍L2����C��H ���Q��K�28��srqұ�?�7��w�(�����^O�wyzqD�{��5Bn.�,���dTۄ���@�a~vo�#8� 6_�Y=sn�#��$��݈�����b����R�˗ySϛoEQ�A��+>%40��G��D�s��_R�zRGq�i:�a��y*�y���BZ����`���>�O��7�N��DY�0#������^H�uD1)��� ����(���c�&���O�l�D'K��c�Ff6��N��`06i�B��9tc�v%�T�EڳyҀX�Ը�F��HO�ހq6�esJ�e,S�����@���mO �#W;0&�?N�ԡm��E0	���.XB�"�o�J�k����.�['|�����of���؝T!�gb'Tc��F�P�6� 4��2s�&��XG/1���[J����nl�� F�5B��.x�آ�"��X!�aǴ� �p�)z7�m�G��	����60n` a$��n_y��wk�	�?&~�L���� ��mĽ�c����)��^�%�F��_�o~W�Ь]�X�����"e����R�O�B��Ms����W�����]�jM�	�p��1��_,���� A� ���3�t���ڞ9�9�_�Ug_u��þvZ[�g��������E7�=�h��9�����r��jpq�imc��̇�!�B��ª��Y!�7�.�5h��=�V��=�L��{Ʀ�9��n`�|k����1|U�1?�'��â�ӈ�0ߓ��˫�oz�h�?_^dn?�/���FN�)Ų��3ڜ�z�����������tz�=A���� ���]���6h{F�S҈nY#:�0*4����uK�핵B/hE�B+�vw���VzY+��V��e��,��|�(��]�	Q�� �RvOPu��s�0E2=e�K<^�� �[\�L�"D�0&�Fa��9�A��#��$���C��9�"0eY�o=6��o���N��̂Y�c��.�$sK�ܾ���D}��A�A�Xl���Y",���XNp��ED�I��_�Ȇ-��I�0�����{r�:�f�@��2<�*<����3<��y��yt2<vk籛�W;������x��ѭ�G7��k?k�U=�l1�����H����4��<~-=~-=~-=~-=~-=~-U=~-&U=^�$�x�n�ߗYiF���FL���)�V���o���7�������ͻ��O��������~n������<š[���8hz�^�f�W���X���4�N�^�fѭ��;��q�^���^��yy�n/�SZ������HE/Oqث����#UEOq�6��������Yt��q}�x[������z����>GO�l3�գH��yJ\�������e����	���eo70+_=�V���C���U��m6�z<q���Zp���k�j�=R�MWU�mɤ��M�5�%�+I;��*^��K�6cU�|B&g7Z�f�^L�n���2^�7�ش��� guJ�5�[�u��g�poho@b� K�$�`�r����@�A�ulC���e�*JJ�R�ɞ���(Դ���Y�����0R�O%���ǖ�"��Ѣ��E+u�1D�i@k���9+�znFO��@�i��͞P�SaT����e6EeÓ��=�-��}9�J�æL�U���g��Z��H]����LQ�!�E�h���\B�ň��P���Z����|K�RB�ƭ�\^�a�����֔���N�..��MtS��(�Q�iGc;ȼ=�D�S��k��I[�j���&s@�R�^��@�� ���hǹ��i�5E�{,@�%p�Y�l30S+ ��o�Nؗ��
�i�j�8��(l[fE�j��5�O�{��x�-�#��ō����sW�IEy�P����3ń���bl^���7�I^���
S0����#� k]����ו��8��LQ���Cp;�G�g�}�E
��sH7�C�<�pT��T�X"��7�$���T�ߤ��Reڜ�T�	[�d����ly�g�?�?6�IK��j�x�/ae1�70�	_�VZ�㻄���	����=��}<.���jpN�>� I�N��4O:e�t�����(-~�]��\q�C�:QHB��+��ո��p��/�!�����C|�����O���@��yS�qV	�Gr�Ql�4��C|"��,���� �{�`�V��>�g�f`�v�(2a����zI�)��4���ER����=rRՐ	��ԙvQ����єl�̻�����9?*�mx�#��N�6?�������g��=��d�cf��������~f=:�Ō���G��:�:��q��J�_�:o�w����l|�s B�#z�����B3>�!q�/�K%��F3͋#�[���G������X�A]��c�q�j�I�\/Sd0I=j]���K ��� X���>����d=E������;���df�ڽ�YLsD��d�##�9&���Ȉv�ɨ�s2����G��'���e�$#��߮���.��&��՝Ъ�Ŕ-�8l��!ԍi{0�#R�&[����S���,�B|��7��"z����WD�ڦё̬�פ�J{�0��O��YHM�VlV�P�)�w�6o;
y�Q���z��̌�[r�]�W��W��^�V��U;�+����m�	��{��"�����M���I��=�wr�%WY��{��o�����i��8�j�Y42��oMW#itW������D#�Io'H��\9a�u���dŐ���5Y	<C�$�K�z����zKOhV^�g������w\,j�@���Ue�6�QP\�h0���K������9���ɇ�zY���cO+<��Ù�}�}������fj]P:F�G\_����_z�l��k���Ų_A*vi��ZB�Vu2=V
ڨ�֨��ۊl;+�-�����\Q��W������@���NL�o�)F��������I1�+���	�{[�G�D7�Hv-���.�BW�II�����^L'|�j?f��أR�ۣ���[�;�_�Ι>���������T ���/p)��e�ˑ ��!�PP���_�y��E�����@>|��3��\J��F��	*�is�tI	@�@/�� ����}d�)��O�їY|�L�����#cJW����'I�!6���bUI\���u%[�IN9���'*��`�m���Q��[��HT��%�8��� 9�,�(�7U�$@�}�_B�TZ��O;���!��g883�.NOC�
�~G���xr~rه�7�����v�v��r ��.�O�>E�<���ë�����J�O�a�Y�J���H���>�g�[�lZ�<:��O�k�VZ2�GO[� �m��y�Mp!�,�{}ᶗ�=p\�ZJ\1���[2�\XU�>�crZr�"r8��&?���K-����"�0�.l�ﵰ/ҠN��Ks�+�%�z ]�(.�(p����}	�sq�1�^.�Zس��_�r-���/�͒|S?\���0u�+l�5���l-g��Z��Wh���al��`�T _-f����aԧ:=��ʛ�nKV�j�q�9Rf���ٓ%m�����;q,����	�S!�vJ,>�IJ�x�9���l�JF4�͈�j����;tXʣa�87ϹiùI��-)�(�1�e�����U�;� �W�zI���1��� ���z� �-��V�K}� ��e5R�� �=�x�6�	�cH�x�/�z6�k�V�5�_�x�9����fִ�����Z������J��5�zF+�M*��c6ˆ��_Υ҈-%��g�۪(g[
�����?m�%v.:��ُJ�:d���!>���3a��I��^I&4�?1�K����Ua=K��c���1]�&���k��S��iKmt�o�>/�UL� ����-������+m�X˪\=����V�����o�$�S&?�[���n�4�K�IAz�9��ç�{���[9�md�PoW��K%?�6Ŧ���k����R�P�{��f�W�J��r��%͟�PK�bE���&�����z�l��ݚ���&i<��J���9����9=�'3�Rg6�쾊�!�ﮑ&s��S>��%���J�5�zV��K�M���l�)϶ϕ�����X�(���ƿ*5=W0��;�8�������8�w,`���s��_ǟ��z�U���:��Wq|�X�N���)Jq��F��G��ĺ�.�U$FE{	����Q~�G�a~=�7³>, ��C�����<�#Oz�G�v��ˬ��(�� �48�Զ#��S��H�*H�*HF)R��3�s��z�Ŏ��4�ܘ�����h-8<U��n�<@�*�^�HƐVY|��?��o͂�ij�����}o�r0�[%c�p�=§D!�v��3�IY�Zt����5�1J�(��L/EX��9<�8�}��@�R� ��K@_��Q���X�-qV���O�y�d�{�i��4�G[&��@2��MN���m7�i �������w0�1�
�'���H
��ދ5H�;���qB/��k:��bz��#���4B�4�}k����2�'��2��9|��bM���7"�����\�&U+�b�J:*�����FV5�,~��"g�U�H��J���5eĨ�*��%�(�f�_�Q�ψ2�+�I�\-Z-j�6��L-�&��M=��F�h�z�kы�Q��ez�7�>66��\1F-�16��L1�&�wR�A�Q1��a��Kò��M�u¬���$�G��5	!c9B����)Af�-���Ŷ_�*K)ъI̶�����{�˶����xI�J± �M|e`�M�	���<��Օ�pf�h��v��ZO2��bO�p*�`�}�v���Ujj�l:�92)�j6t	���.x�G;4�<�f6�t�[;��|�*�����/��i|��Z���#��<=;�����G�@vȠ��߲̾�ɬ)�c������YC	]�o��Jz���	`8���U�3��e�n����y���E�M|�lUAR�jU�zz��J�Xq���P�u�X��	�NW�I%-�f�59�&��VT[z�#�O�����:�m�*��:�,����?�=]���ج�qe��7�K<�٢~e�N�r'��
�fq1*d�{��
��V�_��Z+���bh�_
�<��T��#�	��������v�g�]�s���^�J7���g�	�1����~��:�G�{ a򗍻��ᝤ�.Ig@�`б�O�#��\�+���e�����@�T{Ly��"��!�e�m�ñ�
�i��?��y�+�$�%PY�b�s��K���&%<L��U�H*�@����
{)P������<�������"��sP�� �cA�{aQ&P���SCz�'���x�~<�<��;����?d?�@�r�e��f�����9/I���Z���]^��_�V���z���Z��n�b�J�V(�[���b�Z���j��i�`�D��2�7�n�����UՊn��ܔ0^��F��|�Vl��R�e
m�*�Y�6
Jl*G���k�/�Y��f]�,QVS������T7��r��iV(��[Z��M�AUD���2=�5�Aߘ�b=�Ѓ�hfmE�e�0jP��1EŊ06�e��ڊH�cj*���4����b�/���)&���'�P�+F�7����J
h��"�{iO�'s`��˴3�ͤ��X�RL+a��+�8��<##Ni�x�y�=�P��~t�0 �tJ�?> k�Vn�U�Ɗ�1u�ϟl6��z��d�t;���<<�a�z�_4�.~1����E.%�9G7r���k�����aG��b�nHI�vI[)�S��H}T����<�(j�a=R#p�֝5��f��Ζ�ȨMs����L�h�������J"	��)m�7R���Օo�ma�I�nD�<}od��a{|��Tٗ�R��z^�`��j����$�ʭ�Z�b���ńwL/�$�(�)5�P�����š�s�����jD*�db踹֔�%ʭ��\<2��h���0sk[w��,����������t��tld���&[G럞^\���G�N��K��)@���$�ȌPD򵼁L���=�H�j�^�(K�li���UТr�@9Ќ|t��Ρ�h�A�YS;�\�S3H�h+��EAx\b4-�����DK+h%ZRA?�yJ\';������l�̺S���<5ә��	kf@w���/�M�xق�I`�	<�����'�yC5+xr�w��z� ��аơsoÀ��.)b���<����lh��S� �ɀ�7�-D�Ԃ`h�F�Op�Oi<e��&]�@���S�^�iJ9��PV��zH>m�D��/����Ѫ��nso�J����uUY+ΰ�)QR$dC�����1S��|C��%{��[dPv40o����*���D��a�ax������ꤡ�e���Y�`K��,�yFִ2��x�j@I�PDIfK�iI���擯,�I�㥐�Y��aW"ҽ�lg����fҟ"X�g�nٔ��
+�ϊN�<+A�JV��'�W:n�c�����-�-͡=�V�ԋY��/�"���6��w��?���9,����ŗ+�-��y.�pZBGG��v�䳝�08�V#5u+]?�Jo��cƤVw��w�R,�bz`�*3�Қ�x��Z5��
[�I��;<]��{[�Ej&���KsMk6��_�2��ހ?8~c���g�������j�;+ ���h���������i>�F�W�.��A*p𗝗ǋ9���\T�Z�h��\��g��l1��3���w������I3B�B��'�0��p����l%ԧ���� >��|��S��7�qm�fA��G��8(|b�=�^³�-$��r��F���!��,7܀Jq
���Ђ��A��%%_�4���"���=���QX���t � �:��Zb�/n�ڮ��ԁ��j�(��ɗ��c�H���h�f��r�b>�sKV�?���եe���L"s}qy\�6#E&���.�#|���M-P8*I�MF|q2/�_�$-@ZwVA�2���O�SA�F"|^8�&oZv�iuҏ�� 0�2(d#*<��|�tSD1���a���肧S����""�Q"LW~,�QAd�QY�+^�ʀ˕ScP�>���"V܃�vl=5�yT��#���dƦ7��|(��bj���]��L5%5L^�)1�V���4)�$�r�^�=L����K��Ld�l�44��C����s��r��ӎ��@J_�T�ER0ozX��(�4��'�I�N=�(������������_�.�S�a쵊������Ti�H�D-�g:5?�,���[��Rab{�ɴxX2S�.�Q֩8�h������Ė�c���r���Vf�Yd���4����� � 9�XlxV37EB    f16f    1c0dx��]�s�Ȳ���BŇ���l/8d9Uv��!�����uJ��J�|$������=橗�����i���ݿ���Q�Gvd[��,�.��s^��;���g�Ϲ�fX���q4�Y���s����c�tZҚ����BQ�-K��۞�3���7���޸S������"
�+�r˖s�rr�#�s���0޾3�w�s���5�����"<J���:aHh"�+]m�=�u��XS߻���HI���)޺�v��|Ѳ.��3����5"��m������?�i�g�ΝC?����I����1.G�Oǟ�ο�2�а��~hyv��_`{7�A({����#�f��	��g�G��DZ+���2'L���ʹq�ڇ�����SǙa�f��~0�[� So8�}5w�Їgvd��s��_�+�ܛ��X������XǤ!3���{��E�OA����G���$CDz���iw�ָ�P>w~:^d��3@���'��I���wcLQ]gv��$J��N�DIa���oz������m���������
�4�?5�?�Y��8��)`)<s�����y~Ę=�nx�^'�����S+�`����5k��n��R��f���d���߻�-�V�D)�"'�&׆=YnWDp��_\��a-]� H����!��I��0~ځK��)e�+k�TEʉ0 �s�)W���{t29��=�\^���6Q�Tr����P1��� '`��)rN�Ӛ���ut8:�xl�G�Hυz����K/�k=����*ExQĕ�&�4b�G�`��ݾs=�L?�kFd�T��>��ѕ��� �kᣏ��s'(oEʕ�`2P�1�i��LW���������3Z���S�:����3!Rn 1�4��`$���y�9�m�;�����^���&����v��4�H|��eQ��Z�n}sH���@�(E�IS��P�B���(!�u��t%��֣U��c�}�?�*K��(k���n|����#$������R]����b	��%�ph^Ƕ����y�� zdͮ��묂x���nVm�V�Բ@V����[�<_�$F���L����
$t��tQ|]/�Wt��_�~0���К&�f�ʍ�vZ�[;� �0��X�)�g"��mҤēl!1,��F"��k��[.��{���9w~��/C�I�ݬ��/7����n�k���Yɂ8�ϔU���Ɇ����k�Pc���"�>З�|�~�xa?�drzL=N2���z�(��5���O[�k��[G��i���j?}�Ή��w;p�z����>j1��$��4�5p�IPm�˒m��7m��3���'K��$e�'���[�����D�@`4����HP&B{�P.�����2"
����{���Hi�-dޖ���@KDVb�!��[��%T@,�������c����~PRס�!�����M��d�Y�͝m�r� ���hn���t��E�z������@�e����%� �/O��s�]v��";�r��˅�[a���z�|�x7��^֜)�dx�(
ܫ%8F_��҇�i��O_�~���1���9��EJ(��O�U�93�hd��:��hlp���t�����P6�񽕒Gdp,�����Occ����?-Q���2����\ٷ+KU?��L�:�r��҄�3���.<�����H����J��4�\"D�,��0���%蝽0Z�Mb3�Q���EK�n���#=$�����!� ��S�\�'g�Z�xPRܖ`HӚ�B�ұ<����_�q�ŭ�jXS˟� �`Z$���`pm����筑쭿}�V��ʼ�*������Oi5o�������sZ�Rj�`I�E;!)�T@��O���k����`�(�j���,�i:���/���n��WW^Rh�P<C{�����L��A�W�i\��ō-�,��(]�c;��(�-�{Ǹ��g+|E����ⴾ&����a�F|L�`��uR�p�&�?��	�.D1dI��֧�*[�7�l�3��{2�+pJ�Гn���z���>�p�)���61�;�I��8 {>(ZalӤ��;c��j��i��͜K�k<i�&�M`ER� ~žS�C�Ѭ� �3xA��
u�u�*�C]�?Tnbz�NLo�'��ʉ�j׸���~�e�zC<ʒZ�jq���4�?鵕TF��#�R �9�V�}���R����`q�:U�R�X6с��`���pf����LO������{��!#���^��!`���#����	pa��Q1�ď�ة�UBF�㐠6w���|)���J�z��T �6�qI]p�'��IH�Nl ����%�]�)�x���R���T�
z�nor��(UJ����딟*Q��tJ�R�K�50�#
�)A��Jœ&X����K��b1�r��#0�q0Ab�G�з�d�������-��	c�Y^]�0�<��@�?�WX
4��V��/m)�3H1��(?�UM���fR,ĝ
�T�.v*�D�x�S����j���i�j�H����y�fO��͞^��^���<H�$�U�_d��ig��-���Y�n�N-wL,�&�q��'�!=wd�1S;��i��g��3��<̳'��̯���Bf>����m��r�N���|�^�H���*�#H	lICx�M��s�&Pb�VpHZ�#�)ctv�-گ�ۯd��jA��E�-4��`��̃���Ѯ�,�@��uE����^��:|�5n%Ǐy���^���	W~I!^|O��h�и���и���Z`��d��Y�#���r�(ƙ����0�g�G�F(��fNpo?��oZ��a��@�h2��lD�"��C��xQ ��0��C'I�0�����r� q����\W���4�%˘�+���NfR�A��k����Ky��dje��k}Ι�����J����,0��|�"���I)���˥� ���C^E}��·/�u�t�*T\�Uu�*g�]��O���M�1$A |�=�d�bl"A��T1�h��P��q���c-TF�sV�w���^l+�z�͏l;o~ԼQő5�N\i�21�Lm%D�DYc:� �]Na�:�<�k��M����׋�]��KA��WP��2����L�r���N��<b��,���t����Spb�2YAZ%���6��k�"}�f) %��Oס���1D��%^1:��t�1�	c�3�$�l��	��ZR$�|\_2��[�/�t�(��e*S	T��'�J��ésB��?���v�����xd���)7fF֗N~�C�&�&�S�A�0t���̟�/�Rm亐6�(V5!:۱�"8�|�w|ڢ�ض06�����r�#H#�� ���Z��l��	k�l)y�g�Y��K�y�;��{%V����7��r��ܝ����\��@i�YF濐U�5�5�:�M�LeU������ ��b�+?)�.��;h��|�M��II 8�oޖiM����A`�ںT`����bّ�>N9�E},:(�`�� ����!;u8c3rM7u�&�fr���֝�b�i#�p�;3��$����TC�`h�x9�m:��Z|�w�N!}�]�4JR�ۂ1Lh��w��$�$k��Ѥ]��f:4�UO_��O�u[�JvH{�U��)M'\4�-���P� ��
����m��#F��ͨ{Δ3��ф���,w_��8Nb�t]�ni�
�e��s�Uփ�)9Q!�3���d_�铉p�K/�r�D���F/*�ᩆ��ՋyK��K�x�Y�+�6������`<ں	�0��M��^�,�r����gWfT�1	udGUiI���S�:˳�;fq�9����!�n����D6��[y���?�H�YS�*�����s�ީPm9+R6�&�x���֜'e���/�(/O� q��$�,�4�9�[��2V���x����:�<au�Z�ƕ��![I+�-X�87�Ұ���Bi���^<2�n�`R[���ܹ�5ٽG��0�i%3�X��r�B^ݶ����K30�h���:++P�~-F��C�py-p��VF�Լ�4|%�URU�b�(9	��W����r�������h~o?��<	�!������![X�đ�@��xS9fHYME�/.���r����v�{�M��R��mO*ij���Ұ�B�&��oC �Y����(����$�G��/���'�+B(�{�z=[��Cp���3����pVe6�� m.�Y
�N.{�Ey���D`�և-��"�/�*?0r�����q�l�廬���ƣ�����EzELu.}������>%��-&����������>?�^]|�_�N��A�-]��}m ��q����-�U��u�K��,�ez�&���zuZ��ܱ=�˂8��ŎOGlmG����+�(�zK���J�1πkw�� ���c&U�P�C�VHlZ��-��9�i��hP�jIϘfI�x�Y=�L�Y���a2��*��I� �̀Ţc���B�)0hҝq_o�����f��X��i@
^����p{i�gmGƝF��9{�p�H��g>�$�����^=N-�c]�_��Ujy@��3��k,�ȢJ.��D��|k A\�
n!w��\6�Y6�d���L.&g��F���>�p|z|>�<��Yg�'ߟ��~_�'����ѱ5"$�ǣ#������Y|=R ,��#���<RMRM��,��������>������8��ۯ������(m�c�hj������Pl��f}|���Ȳ[*�)�6����nڸ^~�ԩ����|T�z�ץ=<�����A;�K�+�Qr��D܇�"4�!�M�<@�JD�fNcW�~t�^C�ײzː�p�NN�li~��稧�o�q�L���J><ဃI�#P�y?�9,_�
|�C����wM+bP���%�����Mvai
4��=� '��` �W��:���ڰ��^�g��+�n�7�-,օ��|A�_WᮂE����@�+�c?�UuM�W���C\�Kc�~h݇?�����:,�Qo�ꐪ�p�M�
�)��f��v�E���$_Ǡ@~���#�n��:���������_������M�@��9�����t��n=�ܗ�sP>U�s ����g��:�P����;�[xi^�V���5��JPk������"��{���,Ǟ��/�e������+�<��O�!Є�B��Xh)Na2�E0L&���C� 1�7�4�i`�6&@�T��*��
�U��9ߟ͛��'l�M#aw�x}�'�XZ9��-�p
����	����w��Ĩ� �S�c�9�/�(ۚv���A���o���V�)SqOf_V͜����Ҁ�p�4ԣ�r���1�BV��*!�l��*�Pt�d?���u~��~��\�������β�W�<,{m��æ����6��B��(���YJ/��fs��ϻ2_M��g�2�G�^��%q��0I�VV�[��m��6x�0x��Bw�eE��a��_�I-�x\�6v�!0��
!����2�uCz\�
�C�ZX��U�a����U����k���ez�/�*f?@&�o1���.)��0��yn#t�w��;���C�c�x�>���q����b?^ :��r�J��S��*��tĝ�n�!���"�-��Y��\E����:ÛsK���>�����>����W��o0���d��|�tw���4�����ȹ�u���T��Z��X�}ω�d)F�Y$��+$��0��W7���1���?�Ԫ�=�/)dn;'�$����f�w�2yCϺ]�&E���N0��=��_h b7Y�?�G>8-�����᭻�[;h�fȬv?7��%�G�����M�s�$/�N}��8ٚ���h#�t;�e�,u;�eh�f^�:jZ��o�s��lJ�bJK���emr�lI.�]\���k'p������ѽ�>eG�%� ����0�:���KzU�=���G��~F>O_���*ͰSfdu��%i�uiu��%i�ui�}sq�U77�*�&�c�d��VA�ԏ�՝���ۧ*�rٍU����I��,r
�:(��
�J.(��}`���Ak���d���M0W�����vuv[��B�����B�~5��J���:��ϯ:���.�N����C� �)��EɓuA�	�[ܢ��(Ƞ�hV�0ȳ�/;�e�ԲS��qe$@Y�ԡ��e�y��I1�d����A�p��w���s��=v7Z͚ga��q��N���������-���ו��d���+��h�34��S�]����줘n��z��a�|M���V޾4:9�@��B���4���U�A9$����� H}�kw�����G�T�iL5+c�N�%c�_��(NZbPJ��~� ���U��Ы�蕏^=*��r�b�E���$�l�k�^��^��ѫW�t�\�ʠ��e6�^1N	��zP�^�^U��U�˄?��ʹR�[��<|Z��&��p�J[TzTT�7�J�ʨ�kp�����uR,�\����A�����hC�R�!9m��4�M{5������� �� �m���e��&�*�Y����|�۠�d7l�6�m��b���rʛY&�]$Yoh��/5��:f ~:�����	߀����@=X�0ޝ�r�}��[�Ͻ�{��s.��4�������[���[���������T��+�ˮ1�L���e:�x���O�g�k���60v��� �M	Pe�j����-�q �:Xch� ��|2 ؆q����l�p��G��:�)k�l�!�O�ۀ��������P��a��8Xcdb�@��|���7�]��6���Lg��T�7X��rL�́S�zcᕺ��,�`���n	�1���,��='Vr�T�F��5MT��u,�kWRQ��3O 3a#��9愈Q�4f+��\Ӳ���E逍[���� �KJ� �[Jܧ>���*}M��g��G��Q�����},�����=�*�\A����ҟT"��m�#r�%������>ܤ�Em�gS�"/
��@4n��R�(���A�� �R��HQ�"W�	���=���2v0�� [�1���?�
�