XlxV37EB    175f     762xڽXmo��ί8J#�@!M�RES������j�Bfƀ����=��ϱg`H!�V�· c���?N��O�ӡ�Q: �e��$�^&��Z����}:��Ο����Ψw6x�r�{I���t�-��F��}���Х�ʯI蔄M��
+Q�N��)�M��j���a+���k�]eJk�H']z�ev8��I��i�v���'yj��ʑ��<%F{���ܚ�*�]���L���c�)=3v)�2��l7�6�V���jZx�r*�W�TZ�T"��4�f�����k�J*�L��KL�`Rύeg��@���֔�B{��B"/v��ׇ�D�ҍ�bn�\"et��b7������K����La���1/�E�+7��8�֠6�C�f�NBq����\�JD��*=���
t�BJ��M�^ӥ񮏀�
�K�H��rG�Rm�c��y	?��y�l�b�Z�yn�����(��`<>7.���>�[`�EX*�d��͟G!���Jf��.�U�B��5no�:WH���/�H�K��'�эM�����J�{���u�,`Q@DR���E�Y�,�p�I���PiL��/f�����OVI�����$BO��oNRP��|Ic!+gF"4k��b�U�ߓ�}���>��ؽ��my1
�4���n��9,F.Q��㞪u���(�͐ɪG�DLXZp!Z��{��|��#���ʫ�t���S��zޫLj������iPIv�I�X�3 ���݇_~�:��y/�8��ŏ��m(�`�G��yr7�~a�`kynpT��or��&gx��o���ܢ�uǏ�}L��������A:أ ����9�/ky�,��9����J,��b·�4ؔA��� ��-95ǔv���rt:�G)����Q*ɾ�|�I�VϪ�Ͼm���?F2�
�_��s��U�}�Q~89���X�+�Y7~��Ñ_�tY��Q�1�.њ�Px5ؓ3wP.)�e>��(䒺\b�S����Éb9��	�*�Y����9�b�@��j �>�1Xh��PM�N�O��Ê�{��QY���3����!Q�S[k)�GG��ͽ�������O�Ѕ)2�#I��siУ�6k�Dȇ4O��:��wK�c���7�ؠw�_]^]���Lތ&��������͓��LM-�4����h�?·���$3s�L����w1�/Y޺w�7�fcӏ�l��c�����Y��_����LB��+�5��Bc�=f7���q���,d �ʪ�,�,�z���
�Ѿ�����զ������)\	������g��_e�(�偨��`��	�Ԛ�R�mo��9a���YH��4����^�����̘�R2�=FR5�j�?(oN�;�~qz��׈��Q��P���,�U�e�����_�0�k:��ű���pKB��TyG�è���԰�����O���|�bwT5)c)���X��ȭ��zM*`*��<�^S�0�w����OJ���P��h�70����"��U��K�ZIғ��o�؟��OeF�CP���d�
����X,�����M��А8d! x��L��I��ջsj2[18�5G�Xst
��^�����ٝ�/"���'�7�����EƎ��$
����J�\�k�� �6�.�E�Z�!ҕ��7ѕ�
ұ�X� P�^G3��k3!�ލ�w�
�S~�\�o.Puu�rU�hJ��2�m���.�I�<���f����}�e�q2b��?ۣ�"/�)?p��;i8�:��Τ�1��ޟà`08B�ۏR��*+�Xj?ʃ�8������ך[�t�����3\mbV���J�e�� ƣ�^��ނ���_d�l�����