XlxV37EB    8fa5    13c2x��=ms۸���+0��DJeG���*%7#[rNS�I%���ӇCI��	M�Hʱ;����|@�E���O��E��ž`��`:�~w92.���l�v���G�0^���]��	�wk.���ݲ�@:��m��_u:��]���NNz���L�7�����U�i��Ù1��Cu+xzez�;+��`��
�ŮS��9�r<ku���m9�-2v�$a`ۄ!�ģ>���yΐ���˦�yO{���`��o�NE:������Z���ķ���l��)r�z��Zx�m��VD�4�6L�zD7�Z�v>��&�s��Yg�3|������cC�gҰ�����d�g��y�|G��c����r��Qx�$���$��[�������A�Xϐ��]�ڠ��( %�5�bw�\.=}S�ڧrS�;�YAS��ʺ2x�*��/ f9+�D�q��3��XY~@ͥ��c��מ� �vo>�xz��Y��5������1�2�g�
�6s�y@#�:~/��\a�rL��ݧ��p�1��v��8���\o������S��O�u7��*(�H)6 ��X�u�g-�P9���R@��Ȓނh-I�ٔ�>}	��J�Mp$ �}����g~&�b�y0T�[�x�~n9&�e�9�B��������f�=��
���Kj�?InP���r�/U� #?�i2�
�1���B]s7�z����Jz[���4w�`D�@��҂j��C}2�9��ܬ��[�`M��<wA}����0y>�N�]���08��TE~3���g��_�ƛ��uqs}���M�m�=�{"��hԯ��Ŀ�`i���Z����CӶ�/M���-1/0G/`<�ar�����a3Tư%`��3W�&yd� �lý����q,ߺ���9�ѩUa`?��.��6=>};��W����k��#�Jʹ14�QK�S�����-��c�˫�q��1�m$’�x��2�Q7B���6�~��f:2���_G�H�xt�����}<}���_gR���w����и\�/?1WP}�^0�AS�-h�<t�� �V����s�vػ&6όb#�]��<��w�s8�$VP>�	s����umj:�daC(6b+�$��$;X�5��A��h��E�փN�!��³�2������=J��b�5�����9���L�|�s!~�Ş�	�C��`���z� �� |-��� liD`�S~6��-eIAD�s	r��JR�1�vJd�c���o���J���4 Ps�T ����t0W�>nC0��B��� C�S�8�6�Ɣ�Z��'㈯��Ԑ�Ĵ)"ԅx͓x?5�H����
�=:'�8�\+Y�AB�<�CO����0���|�Fh�XO�a�y0CL
0��mց
Yx��K����J�/!'Q�"�y�/a����\��3�.�<�"jNO�fZqc��`�c��˭��~�~�xL4Mf��}����/�)�Rߣ%y����R�=�~�^��b�Y`8K���0Ƨ�������ӭ�%�9����&��Yp�`�����s�n"����^4N�K���R����)��O��ͤ� I#\�-P��B2EȆLD���)�0%�$��ÖC��Y��b�OB-g%N��z{�	 4d��hޗލ��3��nr��<���}40q$���!��p�#4i�N�_����zn#��D}>g\F/"���O3~0��'f#|R��|�� �z���(��lҲH ��Iu6�Yo�d+�LG�<����ʏƔ\�(/O����8"<�E4�J���
B��cc�g2f��"r��|��|sT�1HLc��6�9�!�K�Q>�Gې�������'�[@$�,��n>^�pBYZ7�%L���	_�)�^vr^j-]�.r�2�l��񿟜z����y��z�8E�`���J��~T�z�w�8ؘr$��/�',����Ĵ���8��+dU5/���.���%	�h=�UN!]�}X�1j��2�y���)g�'4s-�N�;��Bn7��I�t�uB��,��ēB�&��mP��tZ'��ӳX�ǣ��յ��ínF۰
}�Х�R?>y��,.�Gcep1�2դ�؞Z��8R��/�e*��̪�)L�y%��;�h{�����"�"����5���⎂n�b>S��y�#��f@�myTL���O�l|���z�kb*ep=��"����da�����ڐ졽J�K/(�d��ʶ��[��M���xq���f��f�݀�<��I��ށO�|��N�%/:/�}Z��Z�0FpE҃�)kwʁB�ݬ���|��X&nhXR��{ 6��^N�k)�:�8J��Scxqы�@x��Mn�yy�+���� � ��X�����>>�J��Y��),�X�h�Qd�� �h2�Z�xI�ބ9/�$[��/�N'iFm��o���W.���.��H����ts2���u�$y0��(q�h�sj����1��13�ЗF�j�k?�����O��[<E�u:j�RW3�

i6M�T�w���`X��������_I�}���WgW�*ìN6�����!`e�u�3�*ï�r��|�UZ%_c�|�͵d{��_���wO�������o���w��2�:ݝh�a�i6�j2�~x�v�5���7S�����x\���U�6L�6�4�"|������a�������
6J��\s|�,���������z��)������Z�<n��X��㚢51v��??c2�B�5�,s�k��������v�:��#�� !g7SP�?��{���tia��:�)�k,X���"V9���i�>SӍڂܧИT�C�j��M�0IF+Jym?��"AW���f( Bu(~E��)z('�*c������tH�ܛk�	��c��nכ��X���z��I�[-�����M��~�f[�ZD�����	[����"s�[?B�t�Wx�U�)�h�G�`��>CPA�qҳQ�4�:��I�)"��]��Jh:�a����q�	P�4uĦ��[ۡY�`�Zd�n'W	g[�P�!���i�UT�
�!������Pf��?7���<7䚄���RJ�*�	�E
�Q'IJhl*�
��N�&*E�y�
���sH�0p� 7��
V���m��z�!��F�F��3�J�����P�#c0�M��IX�� 5-/PlhZ�S�J�D�R	 �/&��F�A��qV^��1x8m�-u���4{ 9�V��r�*�T��)k�� Ks9�������h[|��
u��j�	%�U��T�~!'�#���/��nAm�U�ʯ�:ۭ*�i�$e�Hz��`�f�*�x��՘4�pVV:��I��I�O��|Ǔ�}Iybz��7��������G׶�0~([ú��v�`��՜c�N~���,�F��_��|2�rBz�B�٢s��x�C��Z�[���RU���&9 ϱ�����'���:�F��_�%��iD����tH�!Ow�X��t�.)f�;�<-=�x'Y���t�ɗf�Pʳ��@�U��ti�=r��Q�\����smE�XsNp��A1���� ���"}�-�ї$���I:!.�2�$�&��z�]�$SQ��y竖�J��.ͯ\bɮ5�#!�����|������8��.�B	�=�E�3�3M��%G~X��âK��Q�Y� �K4�"��v#�]{l5��N�����VctW��&[iv�u~�M���w䲘�hN� jn��srR�GZ$:(¯˃���e�
�R���,آ��5�n��3?��;iH����~�	&�7��ƒ(�dN��f_hU�<���T�DP���Y����tt����Rڌ��lKF�
���Ȏۙ�4��%��A��E�DiR�5��fᴶ��,��4<K'H-L}���a��4{��L��ɪ����_E�#��J
А�����m��k��X��_@;/x�������ɼ&?��2����V��"���އ��!~7w�?�OONO�}�/�5�z��j֪2���{�y���3�cy����S�Y�Z�M�����2n�[�ҥ�cK��&���A��	˕<�o���3��[��HhR�MW�J_�`�-G�v�Fr�Z^@Fi.���̰<:����\��C���eB�}d��D��C�P���>B�G��}��#�}������>B�G������N���c4��S��c^�+�2=~�I��^؊l�t�4�B)���%^΅�G�_�r��Z��N|��
��W�1m����Mh��	W�1��k.Rr��|R7:V��VM�O�Vc��kS8���[�G��I7�E��4�"r�b�&_ǆ�F�R�Q��4��D��-j4�޾Ut�CM`a����;7��K��2�^b�L`e�B�-�ß�
<���_J�#q�ٱ�2g��xt�WqP%^P�w�ˇ��)�#�e��a�d��,�<�q7���������_�Y� g�����	c��Rz�L�z��;�@�Īl���;葅�|��D!#/
�f|-���	����O�*���E�	��t~P�D�Lj���e�c��}��(7SP8�����~�U��W��)]�5�]*�x�n�ڟSߟS�/<���Զ���-�� ��s��J�l�V2���ǶR�_��R���
���Z݉yX��z�PyWI��T�y�8�ǝ��R���F:s����� qg2�o1Q����V'������֢�T�ZT��[P�p�*:z�>)�������F��ڠ�>�Ei��lJ�Sͨ���l*<L��4���-�C���l4��������Cjϛ���L<��J|ܟ�ӝz�a�oS����0E RJq�Ga����F���e6�w�+�:��"�V����gy���GlўRF5�+G���؅� R�P��c���9&"_
d���q�'���bD�o�,�yVvvrl_r\�������N�~��x���;K�}%k����,il�dv����p��z�?�����