XlxV37EB    ad60    1e13x��=�s۸���W�;��uZ�I�ݸݙ$v��M������͎F��X���r��� II�/IN�޼��# � H����~�vwُ����W����I�y/:��n�z��l�a��Ag�����I0g���qk����I� r�o|~*�8 �q���D7Ӕ�͢�C����p8�1�dI���p�yI�`�I4��]x��@�z�r�D�4�碌�r|��}�tw��I�L�,>x���&���j��N�A�ֆ'��p�N�䠨��|3�e�*��X<���#gi�����[��Q��}�L���h����m��v<�r%˔}
�nC-?����}8G�X���it�Y��-��y0[0�g�'��C�g���@@�g��-�ǟD�?d�x�. �XZp
�����	�a��@���[A�����ᄥ_�������e
�gw�x
�l>��с�gK'�x�$ (��)�8�����R�J�p�\D�p��'��PG��Y�UA���
Ws,Y%�����']-�4]��2`$4$�EXf�����ūt�J�"NR
�M���Ch�\� e([ g������pɮ�ss�%J���b&�`lI<�˰
#�q1<?�F�h�� ZV8��Au������?�_��������On*f�U$_٠��w���_/��ğ�7������/�٬�������j�w�����H����?��ꢗ�3e�h�ү0��H���V��Yc�t������J�w�����ho�I峻���������\|,�ڦE?����lt9�.zq��B)�(zvx:������/.�g#G���~q|��e]E�/����#R�E@o���O�?���E��J���N�����2�������͏�)d>:}$�����R-��}8��h�4f{^���n�϶��������;�m�C<��o�E�x�{"^\�_3��?9�08����E����1�$����u�Zdb�d%�ٙ��=��
�Y�/����}?8��Up<oB��m~�����d�=���?��O���G�����eޫ�3��=��QX�ߘ�/�?�Cs�&��B#��^��<^f�qy<�ʹ�� H��X��s����0���sRQ���lh����Q��o�T$���t��N�4��Z_�J�e�%2��}g/��xs�wu��xa�	
�0�������UG ���G��n��|�fq��J,���w�pf���M�!`��E� �=?�5T�,��*>����\�o+�𝗈!�d��d���S0�&��6��_�X`|���I���5R�9H�Ԡ�\-���&�����.U8��4} n��")G�V>V����o�/<8[)�>(�B�-�$L�S��X8��]��"zL��p2I֗��\�C��W��}Oa��[�u賅-*~�_Ƣ7k��j] ���_bQ�e���F�v3��q���� ����"]�`>a�G��\��(�F z:̗n��P���*J�i�?�IǦ�n)�X{�'�~�YT�����,}s��xi��Z������q�������<M��N��0���ě�V6~� :����L6�[ͣet'�nⷘ��\׼r��ù�D��]����=�!|��u�|��Eg��[�t�P\L�� q��^[��F<7���>!d��<�y2�8N�E�kА0�u�G���#��&~c��
{�Vd/���`�;P\�E��.s��Po�{u
u�
����k�[U��ѐ-z�����&i��=w����U��(u��
{�U�v�����w�e=�[S��S#�E���J�ԭJ��)�^��>U�\�N� \���wA
��Z��qt�'W"oE�Nz�Q?S�e
��rӈ\u�2f��Pa�D���L>ovݘx�4��� 
����q�����%i���s���.�6��t]vɶ�f��ֿ��5�s�Y���d}�i0���_�n�f9�2 ~�0�)�`�W�m'ԡ�~�q��s���V'/��H���
c׫9�Iq������:V�`:��-�/b�XG��]<�@��Ug&Y"��'��Я��W���:c�^�TLD`bg�^��+t���>�����p�0ׇZl�Ʌ�WHV~�����#+$�[�ꪵ����� 6k����g��&s��_��8>.����8OC��HtyZ%A����2p
����L`~>����
j��J�&��p��ڤM�ߌ>�ߌ(���QpNF�K#_���y���^k��>X����}�XU�1��!OY��-���9zn�=_��� �s{��2�J�|�]e��&q�R`Q΄?
�$�UË��	�#��zP	|I4Q�ȡ\r*AQD-zj9�07j8̎�W����(3[�:v+�;T�;yg��{�N�3�l+��h���E����i�'L�)�����b,�Q�jF/w,��Kdoǌ�e.Y<�}�v�{\�^*YO�� m)��]6�dF[�g|�F����Y���p	A*�W֐A�&���i��4L�r�~DW]@��Ri /[��W���k�^��k�z�_?��/�u�_G�u�_=�����3���I$�g�D6<�Z���ie�bix� l�|R�|���3��t�O�yR����"�>��K8�]<a���W珊�/�+ �1�*\k �f�"~��<�"..��n-�5hU�q0�W��2�̂�R�9GR#T�<G%�#tڈ�>w(�����߷���^o
ȼ�{��^�7B>����n�׶�q�b?��A���`k�lͰ�g�L�"�W N(Y�*�crj[�L�̶Ă8K'��Q��%//{��(��"�x�NI)���Hw)9�趎V)�d^fq�J�|����.�Rw��_�[���;LR
R�4_K�_Z��JKQ:�:ß6���Fw�B$$���N��OV�9�6u���Ix��Ey%�E>4�(JY[.�O�lq���v�#�F�|Y�	y���A-�+^��ǘ	��E�W�2�bT����H�0���L5-�� �%�YQ���(�'�҇f%��{]%ܣ�J�}*�%i	{h�����9��v4�ҡ@t!�G2�:�-�H����r"Z��n���:�M�Ŭ$�hOc˲��i7io�����Qz�5�.�^�F侐'?#'��,���>|Ђ�Y�_d��r��"�6���w�*�~	�ɒ}	0"n�/Z������UD�� ����$���U��{,��2u��(U& /�l�U��!O���j�ԗ����Ǹ��1댢�!�"����U��|`����΃�f�^����>5KZ�6e��1�O0)������i���&K��W�kM�/�2��4��`5�k#�j*܎D��*�m$
�k�*����Q�8D�	�A�#�R��W��wUp|�fP^�ς^�vN�͈����)|JPn�D)8� "�q���Zx���>�d��an��u���}�F�b1.Q���=�̋TU�p��)Sn˝��U�(�ZN��4�N�of��s�@�\��a8�/�ʣ&kR(��z6�4v��`��|�����6_�]���.qe���a�)���F��������*���k�5�
I��<g�箍��0�J�q�Q�g�\�mb�K�-�b4�aVH��Yx�s�N���Õ&�r ��}�l���&�ue��!���!�4@��}(��
�h�[K#b�V5qm#ϖ �M�E�U5j�!W4�|�����`���������ef�6�D�U$��~5�ۤ�
	F$��x%�9�e�j$Js�x��`�K���29{���  g\J?)�)E�&��l *�4���/���]�)�l&��6P�k1s�y&&>�L����^�6E:K�
fjKywVg�U��rE��2��0z\��l�'��;�Dޡ��������E�2?�����N�*~�xf6P�t,����Ø���N^�YVUf�y��Z&
	;�r-:�����W��D����W&���@1	@ɐ�X��g�zuA;h�.��W��a]%���n��I��E����a�ߊ�/��^�"^NC����T�SL�#�b��� %f^F��{5��������Nc �$xҤC@aəY�ғ����7��SMZ	�f9%��n�kU��D�z[)hyo+-�m堥����������RPgo{>�����2O5�J���%���a�@�mBf˨���-���$���Aۜ/.��X���|���5B�łn��&�Wܳ�{�k����׾g�{k�}�^��W�5���^��7������ׯ��X\XO�x�y�m�R��N���^�O�*r�W׋�@'%s��8���3����� �l�b�`\����B����r�e[[f�H�<�C�bt���f�.?U��=����	
K��<��Z�l��u�w�o��W3�3��6�Uj�(���eJ�����RA�����/�l"d���/P�[\�?o|������m-p���y��6��y��$ �݅�eYw���S���8�"/lqK1P0M�y�Z�#��<�^Xx�j���"�V{�{�[i���'4�c��E���š�P����b�̢�!t!�β|��S��R�ª*R@�#��tĒvQ�
Hr���p���8k��%
QI��za��r�eR����
��yk9�����D
Ɉ�W��L�t��,�'����J����T������Ӭ�Ki�.��n��"��e)���o鴭�)H�<�Jg�z����|[����l�L1��K�h���5��]5�SLQӬ	�1R]5y'��Uj��2~��L�ݘg���m�"wD���° ��3���ʞ�Β42
���S��@Ub٪j�t����p�T���#_���g��l�D�_y�+2���[���94��3[�c����o%���Ԅ9Ɓ��e��ȼ�"����A��#��G�M^�C�vw�C��$I�ԳzT�"�\�Ź#�ӷM�7����?b��r��"�1%�Sk?o�n������%����d|��ǩ�A& �흜����'H�{3�K+`z���ߪ�f�\(��ɇ�l\����I��:ߛ��C`f�����D��Q�b`-w�+!�<�C���4mV�N&�k��ږW��Y���n<}��5��I3�Yl6�ר�^�{ǜ�0�2Oq�x�$-|�a�V_�n�j���
��Z-��������)����k�5����?��aF�T|���ܾB%������bJ��h�Z�>�W�܆p�OZO��d��0w�\݁W;R�����,��9�����ty���o��&jevG%O�Z�3cA�,/�mK״�Qz1�e�O�R��� ��4��9�x�4��O��߱m����1:�[&2cN�~I����U;��<'W�8�Z��=����QL��In��(��Tx���x˦c�hrˢ����v�"�(�Rw����:=ue��c�A�J�LL��nڲ�H��,;��"�"ӛ+�XY����H0�T�ÿ�����ʵ.e]m�n�"^�_�䓝�>L4��e���ca���;��6��
��-�&W�b0Qt��&MT�:����<��M��6����P\�/vz�k�*�voH�&\!����=Ga�� ��.ߧ�U��?_]�$1����i��f
��&���M�9�۶�=���?ҁ]G������6\�8��SE)��S��eo��O�>�m���k���I�Uqbl�,p�dƔ�^Ey���U��d���^���#��*Y��Murz�^��l�o09�&9(X�wk1Ҟ$`�1k��2DQ\b���L����֡�5����4�S䒋p���BK�nAKפuB�9���L����3M�Mu"%��U��ot_���o4S�$��k��.N@����:z�ч0��(NK���ჼLsN��=ּe�b��\?x�k�\<'�oY6�8��%��劾�Ev�,�<��ϼ�^�w�Һ�]���N}k��X����
��8	��_`�nF�eæ��3j��� T�UP����u�RH���_�=y��:3|�J-�B*� ��=�?� @\A��LR:[7��bn��bByE�߈��U��U�/�拵��-Zʄ�e8��788TּU���x�
>o��Q5j�_�"��`��@ʐv�)�lʦta��7cN5fxV�v�ݓor@�F�KW�d��X�g���ZQ9��������xj0�Z(��npK�#��BY|��DN��`5K���J9s��\�%�r�=�Y`0{�������Gw03��\�깖~F���*8���hx��s$�쑱����U\��Ϟr9�|��ȶ���{�o��l���<Rvw5(πz]�u��eֵ_	�YڵWʬ�Sei�Wʬ�]U�{��͊.��Ǥ��iWH���hn�����ܿb0[�7ɿg3b>��a�~��k ��/���T\�Xy\~�-��������-q;lۧ��y� �:�:w��3ԋӰ= F���D8!Cj{���GAm�4����<u��_y�B�����wkK�Z���\�(vV�+h�Ŏ��[�v�"�o����`��_��W�)�]��O���,�8��S,Pt����U���JH~�N>j�*E�Mك�ڡ��-�E�z�$�*\�=�I����@��
��;(:;��!N~�u��S��!ܠK��}��-~U��	>��]ro�S� b�k��?g��R{�}�,�@�|��)���'�(��h|��tCӃl�N��#B�lU�ޭ|JN��{�Q��5�r AݷW��i���r؞��]�fC�6����u�ʘ������b��!<�ݔ�C�?|�`�杹=�`�U!D��Zc���'�����j������O	�}�� �hm��/�����*��/���B�*��p����C�2�ۺ���'��o1~�cZ� WQ��sR�t�{�,�)�#r�c���5��l����/�Z�R{���ߙ���x:F�����樄��b��ԏ��Z����r��a�-��1����9����.�fm���u�	�l�$aIϰ��s��e�<��d"�DP^F� 5�p	��=���V>BA�@U�7��N��v3�y�<�E�+*_O�B|0$�H�v��*���%��u�Q�+:n���Sy�ԓ_3�_�lT���E}#.<4�Hr�q�B�8�ߓ���w~�}g�H�,zd��Ȟ���g1����6L����+m�a���HU�|��<�S\�c͜uSUBW6���]��*N2�)�R
����C��k������T��'�>�΄L�'��Oϻ�'n���Q��}��A	j�m�������smY�~v�F��=�]�Z�����vk�#具�r�c��L_�禰N8d�Aemv��� Z����ƃֿ�"xT�����!���-"�Ʈ��_�̍��*$e���weãT�2��a���j]<�ÐO��k�*yyZu��:�~b�y��l(�[�yqp��Ձ����a��hd
���gi(<E�����[w���]�0���L��Pz�u�����c$iC�8y�p�.O��{g
�߷��S̷f[v)na���� �����