XlxV37EB    3f38     ab4x��Z�o����_��G�$�5�"h*�Ar�hr��^���jld��?������N
mϭ?$��ٝ��v�Fc�O��@�=��<��ns���onb�*J���T)j�䤧t��랧�><��o���u54�6���y��ȴ}�?��]����o\�u�`s��9.xrЅ�~v���GSb������D�g�����\�3ݭ�h2�kT:ı\˴���u��I#�5u����zı#N��ME�)�������|����o��/S�[&]}%�#�[w��b�`8�Lk��w7��z|���2� �!T9����[�7GM4!�I��&���=���h"��J���q=?<����ҥ�-��=L�܍�"�����8wl�Y[7|�5��|EYں��P�S=��j$eX��X�K֗j���d�&���8�E��b`Y� �]b��i�kE�\�B;�6���| 6���6�Of�A�A�C��Md�O>���a3/W�ظ.G�(����h���*0�sV����M��s\0�ܘa��gi\��6�ؔsיT��?N��0�d
�������3��A�r6�z㣵uP�#�nsK(S�.>z��,��No��E��9X��	�~�6]C�La5�1L�3w�j��}����Ѯ����u�N�hR���f2�̴�C�Û���o.>�=U"�Xd����q��W �ۿ��^��`Я��触�/4�YCø�n�ՏX�m�g�9=b�Dי[�_��mk���9�}�}uξ��t��w�X����y����{����X�q}fk��_h����AT(�ƛ:������0빎,sI�nm 0u��l�����d0e��?��f;>��](�G	=fr
h�h�@+ԃ� �� ���'T�j5��0�&���]
��.h6�Xx�|�:
��"Ӥ"�,E���]{�>� ID��#�&��k���)ܯ�Ā�;�!J�Mt7�|ג�����r����Z�$L��, yá-t_Gs`/!rs��7�9��"��ABfrw?8='K���:�:��#��P��鈸e�HZ�2e2��iM�]�6J�_��R��lʾ<N/��p��R��X�SQ4V���x#F��'|y�^��#�:=C�L��XVb6*����4-��_CuX���kT��6�}#�U���*R��!�A�:�4�X�ׯH�����%8G�)!qZD���J��w�j�8U��2u��R�b�#��Z"�v�'t[�a��n��5���_}\�=���p\y��C�Q9��B��Y �Q5����ajgE�?���}�px��(�]�}�'�IOl�6�h��2w�4zy���nxs��q[9������s�Ahx3��>'~pDt�iUQ�Cp���!�9<��|��rJ�Vi
Υ�I
ۓ:�!5��{b#�*4f��XXI�t?�:	-"cp9�"p�G'�ب2@�RBF/�H1��'��.9P��#�a~΄G��L{DD\@̰
'\��.s1v$�I�E
�+���.\��+�}G�su�O?�����������
BX�y�җX�]� 4�1C� ��s6�+���F>���*;Y�)��������T�"�+,\�X��h����Q�=���E��r���*/��i�̘i��+�U4h�Fٙ��,�j�ϟo{�mD����.�>��׀1o/5�&�AEֆ j�pC�����5J��@�������O?F=z�E�3.:CoQ�&`�w����E����g���P&>�p��7u��e����[��Q�Wī2�qm�/�K`���d�%g��e��PL���YU���7��@����(�Qu�kݟ���#o�P�(�|�N�a�糩�
�ْQ�]�/D"�����JŢ
�V*�S[��v%,�ڥ*NJ��b*%�_"B�'���v\�d�X�^��]<8͓�#��$�m)��K�C>V��`����7V)�+99�@�L$ä�H4H�E�JT.H�	��J��=H����@��L�ؗX�UhF=�����M�Y�Q��.E ���V9f���H�8,��NIaA�������	���0U'",}a��a��&}������ƥa����7���#vy�jd6ym��dd��CT�.���tQS��`(A��Ŧ�l��H�������q9��z��>HD=���E��f�rL�^&!�d��Eӱ�&�-�������T�!y����v�{л��d��
3��k����v	��߷�fP�݈fJ�{ќœ�h�Ɇ_�*.�*.�*.�j�5�vJ)�)�g'W��.�'���AWx�P��6H���pV��r����8>���?��x�W�_[�B�-u�/����_.��J��b���-��%�k%;9�
�YSs6�@�tC&c�����­a�9�F$I�<%Q��uN��WÅ{��^8{/��g��|/5Me[E�t2�
�B�Kܩ�(ؼ�8�99N�)ɟ��S���rj�Щ�+�*��t2��&2)��=��5|�m�N�m��ۙ��~�9��m���1�>,��l��~�&%���wl�X�[��,�=[j&��@{�2��e�����#,��l�%�:�!_�X`�E����8����Ҍ����9n\��ղǭ�=n���[?��ܿU����h�?����;���q4"� 8�� ��B@(�A��1v�b���@줆�9;�1x�Nj��/Y��O��c��ٜ<����J�
��c