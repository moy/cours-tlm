XlxV37EB    fa00    2a82x��}�r�8��?+{�=�I$'3gמl���pW�4��qvk�EK���Ԓ�c�:�{����7@ �ѻ٪�h4�Fwh4^������Ap���w>�>�?���y�-�E���<>,O����{����m��m���x��O�?��w�fa��6�4AI�������a�x��hQl������ҿ�,�^�y����»�Wq�t����g��Y�<\!��(���h���CR#q��$\G�!P�9��8Mx���~�j�d�Eo
^�7�h�F�+"��ۄY�w��U����*����g�7F|��(���iRd�����$\��]��a"�ŃEl��K�9i@mQ�Y�w��C��Q �J>�y�f��&2maF�_�޽n���q�l$	\w8����֟�W�!L�_F���+�l�ŉ7��ehrzE��Agf��n���r��G�<���*
3o���`��� ې�
�h�c�p'�h�&��c�$?��.��1B�}c�u����1H^�Z�U���@j-V__��������?<��ʠ�� @�A����0MⅫ*��~��m�
B�z'h���Md����d �������$�� ��<˭��,Q���-�z�t}'!�8\9�ҵTqo��RYt����*|VР��?(n���W?.��G],��]E��@h$�Ck�{$�d�-6��ۤHgJ�b��2z�H�Ɖ{�Q-#�ᬔ�Ϝ(�n��[\<xכM�-�<��e�"��
#"c2���:��41@�(B4;C2A�ʿFs�%���������|pUq��o�0{���`pq�&��M^,�Uz/�v���o�5�
��f_��H	C�-�-X���}�j!�U��F� �!o�:�9K����,�_��vF��X����:��xMВ�IMs��	=<YF�qfd�?�ćd>e�q�x|��Z���;����@�s��m�f`v�k�����w��{wv�kZ9L�^��\�s��2dz\Fנ{�1�:��/�j���
5�L?��9����s��`u�*\�����>�
Z��ׂ�v����
�j6��l>u���;b���\�)����A]Ά���u��5����A?����?��P�p�'�q �P�I7�^�$C��zP���o���\������P���D�P�`���f����qmH�M���Kx3L�}�k�vSxȝ\"���%�V
OEН�ճ4ţ+��Vs졃!���l�@�&�,�1��:~�j�L �(\>�{% h�3�hY�f�-P/��'����"�2F�)���;}�ZU�����F%��n��
s0J���}M�2��*Z�H6����UAi��׫��-r� (�����pY��\D��S@)u@���2��Avl�O��P�7w���m~Ww���׳��ߊ̎/�>�&����7��U�	�HK֖�A
�������}�W�[�l�t]l��]`�#��I/�V�}�C�ï�E��S�����Y�x3�Vmd%d13��&S+����M݈���� #\�ٷ0[��A�, ��@�Άq��#�M�{�~W�ȫ���OT<�.g�1@ݬ�s"䡓���$�0˞QW���Va��A��-��Ɔ�3�&�^�YL����������R5o-h=t�? i��A�����S3�~���ؔ8�:?��J���\����&�>A=�B���񓤢�~��+��QZ�H��Oh�mW���>%��PW����s�ńϐ�ȒE��a��Ɯ=Dk��Q�M��*G�4)���VM���8��%ar#�A�C�f�O����CQR�:�	���:S��Ce���һ`�F���|[o�6���p���-5�Ph������7�l�XeN0.���5�:]�y����pew�e�`d��[��nvT�;�;u=o�.��c�lb����H����Efc�_��K��Ƀŕ���E��\
杤`�Y��<����^�άH7Aor]�.��G�z�oc47V���`��I�Ʃ)p�Xb(#�؈����lC�A�eо�e�, �0q���5����+�yU,,��^[	Үȅs'wi��NA\��AgjYk�bI�g��g����e7`��Y��z�k�$Cޜ��5��j݇`�`���\С�>�6/��ͫ�ݠ�G���A�]0Ӳ��`S�Ft�gm�L��L.��4�������d��0��A�aTf�-4p:Ph�0̊ ��#����O�ȮG@���)��A����@'.�rv"d���&8�5�i�4��*����.sQ��g���_Ά�0N��*Wf�@v9��! ���It�²A�>ʻ].��S��+j�0b�Զ ,�v� ���"�x�B��W�`�-t��t�]�L> �)?���r�t���YG�����~�&�_y����yڑ|f;�"���"�m�čX���Vgm��6���n�;�ҁ	@}��:��q�䂸dҙ
;Uq���xź��q���@T������!Dũ��5���\'`r1�����>��F B�����t[U����N����rX ��"m���� ���A�{x=?#���z�#nX��9�u	!��o^�^	L2���$-�!��2�+l녬�7@���KЧw�a�����mn�=�|�{`&���;V�ջ�X"%�{x.���ޫ�U��ܦO���x�+?���%���꽛W�x�̈���<��Ҭ �wʫ���p���,Ԍm ��oz_�!KeH����=k�̪�-��Tbr�g��������{�ǡ�`r�UX�Z3�1�/�Ӂ��Z�B�����Vҷ[o��T *Á;Q[m\�g��.��uy���l�.Og�nü#7��V���3��~�_>�9tC3�E�]SG�\�2����B-���VL��>*��t.�$jK�8&����4�wd����b��;+=AgƨїD��;��r���	��=9��Ѽ��+<_g���!k��)ʳ�=z�;�.sߌ]\��j�ҵoh���{;-L��`�����_m�^�CO��1
�o玵��[�w����F�2N��!Z��*��ޮ��S��p��&��fj^�H���4��a :��cEX��Q��̺@�h�poAW
�|��*�m���Q�d-����&�7�dkR��7#�W�7�u�Q
�$:�,�����o��蕷m���Y=7gr��(;�����(�p��Ʌ^�P�%�~�̦r ��!g#8�b]�%�p���\��<`l��
LlF$��|����f�k&ݣLi�!��	�<t�91���Xܟ��nrkH]��mwJ�gA{س��.WD������C��AfiN�W;OYd>W�O+r�$��7��h�]�N�`č3�H�"��̀H!j��mܰlɠ&u0��s�E�e ��kX�Q3:w�J>6��� N�!�z���)�	#$���g���Ҡ�bAE'��Q1W�`�a>�#�S��_^:�����mכÛii� �f$�)�Wi@�6����Rk��㬚i��Δ��e> `�. ,�΂��W 
�v�^�<%[��1�P(�8�!:#k1�>G5�W�q���lꬊ�V�;�Ԯ��v�. �=A��	��ԉ-&G����!��u�t�Y��guhk-�Ȗ��ZuV�]�_���q�����')Z�
&��m1�h9H
M��4y$�:d�#q�r,o{A'���oE�\�.[A/2e�(���i�Ы��ki�~]P�T�Ha�z�@�fQ�o2H��$�b݃��t@4����M+J�j+7o޻,�d�f_�n�U�n��ؐk�`�W��Z�CN0�ǁ���2UyE�b� 9/��!K��i�骩����F�Pla�/4�n�=�&��7=��Gp��^��'oq�O�����x��NȑC�^G�8,p#E���ՠ�w��Ʌ� 㷣(6o_�7� �`6�t	��.��{�oSQ����f��O[��t��Fz�ҳ��-&�-r�`��6iQ�-�o�
L~Avp���#� 5��x��;�UR]^|\%�Z���hp�,��Zpѓ�yv�0��t-��2�$�~�Ӵ�ŏ�2j�	<��z��(r���;������Edar�4 .�ƀ�Ͷ�R�q�Fq��~�4�{d��7�Y���j��"Pb;F$���2��F�.R�6���Qy:�a��2��ǟ�>��������O��#��?�lҙ�;�w�$S�F��X�J_ n���	q��,I�[\;��m��hsE�����s�J �I,��bk���h�-�TТpBt�"��Fԑ�D��9=5Ԫ>}5�
~�iҚ��Km5����.�Fs�b?��~��l6��٤��s��=Qo�Y�9����\v{,蔋�vt�}I߫��Ԭ��n�u��JҶ	�&ک�
��E��}�1-�BK��H�/j�d�7c��$�	��_M���b�����h߃�þ������ß4�e�:�5�f���x��JWJ�����K74�MΉ,���)�Lk($ƁA�j49'�d��<�2���B��Y<di�ns����&Յ���ꓭ"�t�\�2�$Q�C	z�4\�B^U��<��b�`IV���ȟz��b�&"���)/UԒQJ�_�ʘ�<�^�^�I�at�"�������t>l��k{�h�s�㱞j���u�'C�6������	��14��8J�^�q�{k���q����2�=o�G`��^2&А���#�����JĖ[c,R�8H�A��M
n��Ì�U�_�U#&-�4ej�0� �e�T����	�����0�qb���ղZ����]q����>�^L��w���;�ӯZ�v��z���Z���Bu�����U��oE�߾-�[q_���{�H+�^���>Ķ�������gE�"M9���1�Fjb�y)�!�,�kq�]��6��ߠ��h�:��m�eh����z|���V1�vi"��!(#R�hP=�1|v�YT���{��vD�N[��B��(�n�	�.D���eO�hu.̖v�:�v����R���9�]g��*/N*|\^�
���c2l��Q��lM����ףY��}Q˿\�qy��u�<B��|CW�gV��[������)�)SA.�=7�����i�kH?\��ঌ���}<ێ�)��"Ö����L&�`�ɟ.:Ԙ-���1툾ܘj���i����'�1C+ј�ޒB��`,�6�X}wL�i;��ם��V�`����h*J�|�Њ%�R�wS:Z_��<]�����HΆ��噬��}��VFE�%/Me��]i���"�������jr�(7rJ�XD �fCٗ�>��ቷD��RѤ����̪x:G�b����8 ZL����Q�sH0kO^�Zӎ��z��dH"-����Tk'���?��Ԫ�����ʳy���#D�5KM7顇iZ��Y��XŶO7��3�yT�ŭ���`�J�eie��f6@0���{Q�'Fr"�hF)r�1҇��f�R]�\C�X:r� ʒ0�ے$�C�Э�0�^��t����Sw��1X<*��4pQM(�_�̦�䲿X�ٚb�^Ő��^K����)H����5�eq�Wu���om����"�f�E�4��"1�8�R_����V�"�	�*Ir��@�Dds鋚�#@����}�g3�Sr�:�瀂LGӴ6�p�7�������&�z�M
� �fJc�q������*)�����>�}���+�/�r�c��m�S)#l�-C����Xb��:�����#aG� [�T~�F1��ˁ�:���{�Jc���b(��$���+m����W�Pӽ\��M�M��Pd|aK��2�.���\�OsY7	̐"܈�a�j�ZK*o	Y���Hqil@.�(�&��k9�� <1��60�����
�rFDV��2�6�!��&�,d���I}5E���'��InA������0�tL&��|�H���*�yu3#��*IӣP�|V�|�	H((<���݉�ƛ6�>齽�9G �%��O8"�ED_]ȵd3�?��wv�_م��+M�i��~�b1�����h�ښu�w���C�(4� R/,
��˷��V����O/]�W�I����?��7C���"^����#X�U����7HMF_�w������?�{���$��vSc~����ZKP��.�K�A%Jm�A���є� ��0�di������C��B��'���&���T���,V]��v[��bg��������*x͇�Ʀ��V�|����8�c�3q���rOi.��|H�`X��@��k@��7���!�����o�#�p�~�ß��S,�/?��w<������g���ﮇ"P�֩<��+�������C���w��]$=V-=,`秬L��$&������Jȩ	ݓ���&B!��=�j^~��U�6���ʯX��8iH|Z�b�yT�N�SS�ټ��^�yЛ���-o>�w�~7<q�pI?O/\�>⟧Zk�����@5�|Ƨ5�71PMfCMmV�P~�~�\h�lf��gp�r�^97*�7Xͣ��R�ܽ�v���O:w'Q=�d,�>@�F=/����24Y2��#H9��zI&�א�U�{u'Jt���Y��r���8���@k$	ωՁ�W��ڡ:�l� 7�t<�M�g���"~�xF�Hᯔ���>�Gr%K�dc��n��`�ͣ<H�֚�j�㌷�_D�3.�X�_e�����u������c)4��%!��A J�N��j��$����]����7�>�ܧ�ՕA47��rn�#�|�J�Q٣:C���t���	Sy K�L)��A�7{��Ԃ��;�`�,9�^<g�Q=��_-Z��Nڗ�M�}I�ܜ�Q�J2�%ϒ��W�s�U"[X3�PK�{bĴ�4=p�W�o���r���C+������"pg3�4s� �)�����P�=�i�O,������􀉹�3%�N
 $E��ὑe5,�(���yԅ��h�yE��ZQfa
Q}x@���Xx��)O澡T⋡T℡T+S]1:�����uG�\�r�E�"�s�Ba�PvԴ�+��S�Ԣ,��_D{��v��|u;�[\�  ��n��n[�!~���'.Eu$.>��t�I�*|�/ݺ;�g[��%C��J���q��i�{Xq�DnQI7�0Vۮ&vAh��v�g��u3��va��H �D5�.-�btc�㠻4�yrT�v�٫2|U����U�?�4t��:h�ݧ+~�W�iN	2���#gZ�c9�d��3���Ӣ^����n��K^�(;��n����;7R���U_K�[R����rBމ]h�nPi#�Y���՜��6�A�nE�W�a��1D�y�\�2�2^5�ts��	͊�D^���J��M�u�mB�T�%�Ό���N������U�0R��R�2M!�)���.6��>�:9�n%���	�"!��z���7w��d���O�����u��q�h�;�����]w�tT�h�@�� ׆�ZC�O*�*|?V�Q*���ڕԫ76%�]��ۑTڔw���L�:�*W�٩�}z:�[ ��u�I�[B�c�W`ۓl���6|��A��j&&�������g�u��~#�vU�g���6�O5Q�u�&��Ψ���*�HT�7l�oR&��N����?�1g�z��ս�ѝ��)�W7��a�->�E
Na"e0��YNC�ǻ�UUӱ7HƐ����Mpe-c:��NZ�r��M�з+ٱ5��+P��B���x�K[G��H$��� �O���7����\�8��+h�Ei��������'^,�\K�ޱϒl��my�5��F��%>��^���ߧo�a��h�B��^~�\�1�Cz��+`E�&?PuK���+|i��D11Q'�1��UtW�����A|�&U-
>�m*ѣ"�a��QRԌ|��^g:�\O�qُ��E����m6�1y[�Y�!=9�̅m#��⻂< [���^Tcp+�o�'ϲ�w �}�)~хmV�v���|�/���_��1-xӒ�+c�lK����ߖ1c�1�H���S��#���>�)K�P�Rol{�T@܄�ޤRT����'�͊�I��=�x1���"E��˹В$�b��1'�s��H��
g�K�~S�4���88�qMxJR��E��HE4�@HWCuU��.�k	��b-e��6}��V�X��l,ӥ��2ajyO+�Z��J�ÿ�q�B�>� ����j�A�h3�� q~�n2�X-97���w���r'�����s!�+�����N8�K%����xi��h��~�5����]Jօ�kuPH=���3U0
�g���x�����>�ᒹH�
���CR�#�1��\H� ~� TAhʖ�8��s��#&=�m��������@�S�J�c�L��h {C��"���	���.��ҝ�X�(TN��>k��2�=��J�di�+=�����ÿ�������@�{�����-�x_/M��+���8�Uzc:*�#�@�hH��?������'�)��N����K)��"m;C��;iKQ�ݢ?����5&8Zjֈ�_�V�f�;�+ _����M�~��:����c��!�4A� ��a�X+Sn�e4�������Q�>�ȅp:�gM'*h���������|G˩COJqy�	h��D���#A�|����ީ�#����Z�b�d�{&���}��ŧ]�!`����/��D�������M�����i8$v�÷3�8�D�ȭ��(��Uyޡ~Է�S"�Iв��!=oĥ�6@�hlas2�
�ԷR�V��'��#�?J��x�7��xXC�)�ޝ���c1�fm%�x�g�]u��������*/������}����M�}諆��>���tyn�J���o��l�C&����u�Dx�}���
?���ǜ�f�wwBp�!�$���J�Yw�z^�Tn`�Q���h<G��jґ����~2�/k!d2@cL�O^�S4����@��޵=�'��^��w�\�@��x��0���q� ?��h��I�d,���Sny	M>�F��˷��������*�qPY�P,M�1��'��z4�>��4�G�^���� ��u	Vo��:�S�O��$'i���sǙPFЀ�!5���5�"Ӡ�0�0p�b�(%����$�Z�m7�w���l,�ő��S��ڰ��Ҟ�gP5�L�d���EvڄY��m��j�����ԋ�ǋ�pP�zD�ҤG!.�e���$.h#���|�v����X^��@۠o7���p"��ce�p=��>P��ٖb�A �U>B��2
�)�r@����-��,�U=�Q_����C�z�������*�t���;U���)��MJjXGߎCg��쿣���Vݫۻ�X��U89M�YI�J�O�4��.�E�e9��շ+�}!�"�/���M�ƾ1��j����r�Sl.nR������9��Z֡0�:�����냦��܇:��B<��Pd���@��.�O`���u�'I�B����b�p膯�(���OzW� �tM�Y�W�<+M	U��R����,�/�<�|g��v��Y��^^"y&qj�[s�&�*�V�����\�s�}�?�q���I_tWl��%���H�'Mt�eɋu1O<E�1Jz�a���/�0�byF�Z�b�xI�o�;�~��hýV%!��]/�Q���iBrͪ���BS�V^l�9MU��ҷݳ��¦�gSv�_�wy�"���scך�.�A-�.~җ�G`�//�����60}��N�������S��Z�ea���jW]�+�r�[�h=�8�#f�� � ��#9y`@O���$� �t7�;>;��pa������ݒz���"���;����$Sَ�ozY�#�uu-��Y�GY#�/t�4�f�sK�0�����|�P�}0�W}��h;�j�|�����>k/Qa����xz�}^��Y��J��O'�kB�Ž�Y0���E6�C�Цj�Ze�m��2H��"�͂���au���dA�Ur0�BuӼ�)[-���΍9b��Ȟ ʰG���:,J{v��H7OPm�<��4,���F�}�m�y�9�RT}�n���`��\�*��-"dH���P3�{��Ȩ��S�4�?�1D;���9\�A��q��%:J�I�&��;��O�;=E��'�+~gВZ���ܥ�-{�����r/8�R�x�����U��V��]J؁���/<a�0�o�%�W�]�Ȥ�G�L�Y�6����Ik�_ݐ�6��%�oJu����CzKvTC��'����C�?5Nh�����]�7���:��CR(�����B:�����FA�&)2�aD%ӄ/��H?�|����h���>FxL>I��]y�'��L�A���BKU��&���>�r:<�4����%G�E�Y�8�@n4!)�|'�� �pҫ=���#�QwA�O��0D�x�Q�ƛ�ɂ��}����CM�V��ݭ��C��.B��Y�H�N��� �o"���Npqx�����D'w����)������%��I���7�R���9q�-�RƓ3��HCؑMM�"Tڡ��-���i�p��C*��uq��7�ȵ����N ���F��<��`~5Q�z_���IFXlxV37EB    fa00    220ax��=is�F���+����.�&@)���T� feJ+R���[(�%�)BH[��oz.�	)�����$8���t�fz�᧳N�Ӄ�`0<=�ǝ�
g�-��f����QЛ�Ӡ�<��M4?�h��~���yй`����]�k�M����g��^��i�[��Vo<��1�z���v��& Z�Vt2��3|�K�Q�e����ݽ-�|�r�z��p_�n�ٜ@�G�8���*B�y�ID��cp�ێ	�4!͒4��xϮ��m	-c�AD���7�x?��Y�S�Eb[C�E`��[	�ܴs���
�*��7�t�f��%��.���Ŭ��i|e��N�EQ�X�����8E����Ύ����"�=�h>�4�7��i�~��}4���bʢy�����!��)F���A���0�0{��n�d�,2���p4Ǽ��������ʛ<$�x¤���A� W�QPpwi�������3���|��X��=��=_̌����D(R�!�Q�:~"��Gq��������q4J��`6��t�>gk�i�
l�.�6B��}���}�~F���fQΩ����^�9���	]%�4
g{r����٢\�����NEX��r���� ��ǰd�@�O(���ir���l̣7��(��d<S䀕i���|@���5�x���αx@+�w�xM#�-&!��J� �m4��ۨ��6���$�ԍ�빱���A#�&8�n�_O���ӓ��t�ؓ ��<�^|:��Ó�1z�T��`S�a��ZeC��RϨL��4�c]��l �4��NC!B�(� oy�\��A�H&��ǋ��������'u�y0��WK� �	��B{��3"4~�Ѯ����(��م�64׫��Q���]��a�LX4�_�HY�}>|L�:c�ﹶ�A���@�qiɖ�X�ŝ\C��]Џ�;��J
o���q3�@�V�p�$�-V"00*bز
@e��)�Wa��
��M�(lY�P-s� a�Pē>Jɺ#��]�1t����h�ȧ�V5�����0��J��`Tu�l�Qf�j3Z5��y�$Y�8�I�̕��?椀����Ŋ&��(?�U�rZm�IS̎d��f��hm��t)k2�YS?������hBE����[�lҶ�$'�����v(YK?��C�Y�Q��OE��+�������BL%��"��`��"�X']<��Sc~�_�|:$�^rq���M��ބ,pE�<��(#sD���֮ڊx��I&��=�����'0([��ILA�4��� p���;��*��h.�����y�b�� �*���p�7y�e���=��!N����ˤs9/�����T]����VL�i������� D�x`Y�7ւ&�F
��禉������_�W&Twe�艕�[��
�H��:�{�m��Q�b��z�0G|:�@�i8�Љ�q4�F���&��Q�N�ՊͮM��bxzvtz�Q�t�痗t&��qi�o�e�fڀJc_���!'KP����9��ܝ��%�AEF [��\�{��j"؀�r�$�J0��\?K���Z�ܽ�z�r�k�W�)�u�5�-�����㣜adk��B��T /���؂���4X�V]�W�׶����K����رz���)�޹���i��8eH�&$6�x�\�"�l�z�U�ے����e"��ˁXr�Z2v`�ޚûY#���YxV���y_��
���{�pr�F7������x���Z�"���2^EФ�&��ao��}8]���H�&���z���p�̆�\*g�C|T<�Gi���gm5��W^5�9�gU9,cSn2�x�=�牠��kj,urB���֝�ZB	��m�7j�$f��Y��h���b��(D���۸���b��� �Ph��խrӎ��o���+�g���G���E � ,�ؒZ�B0:�0�V�^�0��s1��a(q�`��i� Қ�3�3��q��G0xɢ��	�u�-m�4"k4v��k�)�gf�'��.#�I��O/���B��Ƙ�i�(	��f�2�΢zc��a:t�-�G+�/ħ�l�8�x�z�ȡ�z�<(�[�L�υ�`�i��g8L��(��9�z�]fغI��7���3K431l�?����bJ�ɹ;�v\i�`yi�4��l�.%�ᔅZ�"8�@<��ɭ��˞c�lՏ�+G�����?6մ�![\�t�r6Dr�ha.Y�.�i*i�1��H/�s!wb���Y��n΁v�y���]'tג�o�o�{��4���rΨ+��1T5V
Gi�ٵ��sz�X��+�]y�8�l�Z2�,9���.�-Y�+\�sgiy�v�~NS�1� %�܇i^�I�8��l���O��Q�ٶ�]n����4�G��1��lo�+pW@(Ӷ������_��_�Lؚ�H��im�_UgRԇ0�{g�{�G�=�!仡��ޢ�y0���fbmqV��x��[���5��B�J�H�r+a�j��	Q�,�Y�Q�K�Rp����
Ն͈�mh��$K�2f��<��C�!�����d6}g�z�L gd�<"f2.|�)�q+T�p�HT���)����T��=� ��� 8���A4�Z��N���䐜;�m*��}8@$��"�R��y�γ��v��׷!z����1H�� �L�SS@]Ã��!�<��GX�s��t7G�@�Ư�y���m�诨���oq:���R�|���P�'�G����Q�>��k�/�w��m�=S�s��3�|�7�}���v��`��N.��aGqi��t�����O~}���S8��_-p& ��=�]B/.�>A��Wx|�i9�0�i�� ��\�Ɖ�r�|��)M%z����p� A�K	����ѧ����AYޯ	߮D>����`{��ŰM�4�N�� ���8栨�C1� *�R�G K���8��qȣH&c5�X"�È*���h�G�Se<��MzK:��M�����T04�x-ã�'V�M�tUNwN$�ݭ�l����Y�;Q�tH�n���Mw����3�S��"Z���sخ�a���m�i����N�<!^ey��_ޭ��nUf������\�����wu�|G����Mm>`�֫�r�O�_sXR˹�&./�gk|�Ji�%������si2yyz~��z�l������O�?�x�#Jvn��f�R�, _�Q��9�����{o�h ֻ�̟0��ZYz_ê�⫧({e���{d���_�9c~���^X߀Ղ �5VKd�ÝW{�pV�^��Vk	��J"C��-���
w��ĺB1�%V^�v*����v_���0�,������X�����L��w�n���V��
���BΣ,�&�C���Ekch�����A��AU{x_d�:�j�L@a
��.[�*d�*p�p��4�����믮^u��+�ׯ�^��z�:�������CL�Ax�B~J3�\�v�f����_�@��~9}�@�h�F͜��$��n��b2��t��29$��o=�Q�(1Kf��m��Y�e�-�u�b�t�n�;�-b�q������yD{ΟH0�zfy��Sh S���ft[X����S.Ŧ7�͈�1#�=�9�jFI�+C�1`*"���T�<���:��r�`����GtGvw(�J�#����cz ��J$�p4��L(e���tD��
��@(�2�J�aĩ�/�}�݀}�,�&l�a)z�Z֯[�FՖ8:ica��qiިNȐ�Z[�>��e��_��w���]y~�/�����G�c�FJ�O�,JqT���l[�dޯԟ�κի��]D|�^˜�C��Fm�Gh-��i��I<��^�K�%���m=�^6�Ɣ_����)��-��T��6���!��
]�Ǥ��ς;���n䛹�d56��/���oН|���u��÷.v�����p�=\�T�`�0��):��/lj�yr�Jx�I������Pz��%����av~��B�5�����\*�����5=�$>�߶L��2��C�T����h3J�\��I%a�ٓ\�i����6I�0�x���(M��"�k��;������8�Z\���%E.C(�@_�O���]F�ؠ<�VKfd`h���@9n�����8�$��,�n�h}��io2�����P�::���(��w���&Ỹ��u�S��k[�z�V՝��c"9]A�8�&����P�����Q����h�&�,"5^"vr��݀3
X���+��aA��|q�_,���p#�����tf<��f;yES�f�r�ڪ]���^UFF| �`gM֎`=����̤,)~�5��mX���l�~�j��E�%��a�dA��}�Q�7k����Ȫ��.��R:���Ҧ{�W����b��~b��k��ڞR9]t��B'��=%!�}IGL�<���p���M��7������+%��/����Ψ�� �R�`�Č`�4�w�� k1�e�m��+/a��+�扰�NKDȝ���zP�;.�����慽h�z^�����5W6��vV��P=k�����a���-}���|t�]Ct��f���z��m-�{p�������rp6c�k�׹�ĭ	mʱu��*�(R��������_=��@a=����B�P)�b����g��4�̑5X驍��,<0��S+s%��,��	��J�*���+j�oo)v�m	q�e�a}-��G�����.��t�v6���
�㫷Rm+^���2�κ��<G�p1����	�`u]{(�5c��ώ�7�m��u_¢�Sؒ��+�"�k��G�C2���Ej,FVj��gl�{t�>�kXb1H{�z�B�Y����m%1V�-;�H¯���/Ͱ�+{�V���P�H�CA0t9�+�o9PIU�����0k��.�5(�:�u����[�#�C�
�U�SK��Ep.n_�Cg���W(�ǎ���������V��.�Gg���%uk9$%���;O��ɡF��ے챴;'�Q�5���hʝ�o���ќ[�zU@}�]�������}����������g����䯮�v-5����e�Ta"[IM~E5������}����@�;Մ��nB�M�J��b�W(��X(l�u�[��8�ϟ���� '�ȭ$����x���my�]�+E�\Xe���3'v4%p,9I��+޶����wl����6p.؅VX���ޡ\��
h!�4�7Z�`�]ơ�J���l��#M��k"w	ߒ>�3�*A�_		��m���m���U���e�j}y����n{��Y�v�5i�]W��J�}o��kj���]ͭ�T0�B��r�����k�u�R��n�Z���r�}�^˹��jUm��ZHJ��(_b��[>��eV?@f�jfV+�ŗӫ�%�Fv����P%?Z0�س$���xgA�W"�C�" �G[�U+㲥O�W�>��I�~XG���(}���_O��n�}�_�>�_E��%}�[��'���˦O���'=铿��ɯ�>�z��K铈�������A?���Ҽ��{���g2�Ά���RQ���0�>5,���)=�%��ۑo���x��p��:8��P_pI�y�[�W�9��t�N�*	b;+���Ypvr1��,��~�i3vO�8���U| �G�J,��=A'��3�8�Ήb*��/�e0�aFܵt����m4�n�4o�����f�P�t?8>\�k�	"�3a/��j�����i���H���_KW���y���b���e�,k���P���U	_e�v��i2i�	�ȭ���߳��~� �r����_��6�b�*.�T)pw������`d�^[A��| �݁�$�0ڏ������i4�7��9prB��Qǲ��<�� >�b����N+�߀�A���.�u����ʨ����!�_A+)�H#��Vx�+I�cX�E�X� mo���X���%׎��U'd��)6��G�n��!����{��A�	�����9,��w�m��%��cٯ�A'�]o<Q=B�F/��
��G�#87n�J�����$� ���&��K�NsV}Qk��]�c�3/�*�E\��Y��PAK�Gݏ�ls9(��,	ܲ�Ds�l��\, �EѠ�MiE	~��w�\�Ri$c\w�pN7XË�]�JՀ��xt�GD��[l���C�DR�@AKS$�+Q�D�2�.�g^m�Tn�]��tT��uҥ�xb���ٺt�:�m��K�ɌZ7�*����bx?�inX��׌O�3����j�m�!��>��2kN�~]_I�!��2����Ь�84��sW�\�̭�:\�C�Vez��E9���K��鍧��8��ZfA�B��&�����I:zB����&���>�q����9�2lx.�)!�|���
p����e��yo[M�#����<Jo�YD�����֘�b�g7�b:F�YD��(��8���(巿iLhTԒ'HH韧ZpK�g�g��^�E�*`K�\�osH�`�倓�9���P9` ���$	1��h�aW�c�$J!����R��!�������J��
OHBЅ;|�ܾ��_,���]!Ŀ`-�j���޶��O��;���n�R�7i!/��}��_�,��K�@�;-�WQ�Vy��7��/��@T>Wr������rH��� ]jQ ��<Tʊ�8X����Qp�ѷ9}x��{&���Q�À��{W�uq�k>z���i�_J�Ö��Q�RP��]�)�m)!K��{c~���{t�Q�b�#�>�2��ƨ�1x_T���6���G/F�'3�W�C�S�8�M)�N :Ǐp
/�߸�$W��������y� �D�z�)����5�6AU?��R#O�?�1?��� O���S�#�� ����?,)ڛ"t��0�;uq��ɰ[+7p0d[_������h�VאPɏ%�\�4,��i�����0,����U�#8h?�g��W}D�L����?�o��y���C��A�~+F�Z�E�F"��i,(~�x|n����S������2��RlyY��c���+Ny��!d�4Y��N� Q���<�9�
�`�\$��pʟj�f�4��,+jD��Z��	�bF�V��E����+�4-�(�Uyf̪���*���XZf����ϊ��>׉�{�Cp���G:�[kQfv�"����%�����Sa�D�A'E�x������Q��8�,."ˁb��p�Զ�Ӝ
��b*��T��W1v�p|KS�Q�Ń�M������N�P��?ῠ��C��+�2������﷚�c��X�*����Mng-�Ǟ�����w$��hZ�W	M�}?4�C:��<��;�x�����D�*���;���S�k٥Fq=�G��P��bU�,�f�\�c�ﱍ���b�}�����v�K\���m�U&��ek���Z�k&G��r|����E�Fc��*���'F�,�����"�`A���J[��d�'"�� �6��}�X���o� ]����h������
k���[_�e����=ѹL�F�gP�o[�P����'��x\�żf%:!a}7!Q.7lp҆!�/;��|�ge+�.4s��)�2�.{`h��~�L�%�υ��^��X̪���0.��!�U��'��W��dX�g5ǒ�M�[��d+_&SbȂ[c�s5��������*)���5s�9�4���lYٵ��
�Un�z�Z�ϒ��y�i�E|�>U3��n1��۶�Uk�&_�2����e� ��8 @��%�ϥ̈_獒4G��)Ȧ�< i���r�L�L��7L�+"vɸ�k2�M����F�Q���ujm�1�72��*�"�[��?��a�j����ò�:�ꉚ:�i���ᮤY�_z��a3,ӵ�У�C����B��W��CWl�s}��m	��lw�����d����.��ly�b�U�.�����X4���w����
5�c�ҷ憍]]�_U��&�_�p!]mnV�Z��=f�d�/I�oC����7+8����W�]��~��o_�m��ˢ���d��yh�(�(��YFM�R ��2�����	�KcGA�7�x��"���W�ʘ��c�N����X�z�H�T措�u�P%��,�*敂�J�%ü>�;p������j�KY,�iS�]��q�rޤX��/Q$�2���Y��BQ��nR45���~�)1eK�L�Q����T�[��OA��|X�kYE��u\� �2��aT�I��lJE%]��~ܛ�?��=���EBV��e�|�ie>e	��s����r�u�$p�7]��WO�7(j�=�|v$u��0�}�(�� ��L�+��6"�o���Y�k�HhV4�\8ͪ�J��9j���V�VQ�*b��I%�����p��+_�zXM�mS����*!� h=��&"��~��xF��U�[��;�@ghP�ri���4������쭋e�����d�b�jqG~N�'R�LN�i]���u{�1(1P!h�W���7���m���~i�%ҚU��+��Wd�]�}�$`����Rv�7#6���v�o̹���zՖ-�Ǽ��~1j�e���yp����� ��4XlxV37EB    8c4d    1566x��=�r㶒��
�y���wD��V�N�m�%��#�s&٤X�Y<#�Iٞ-�v�F )J�&3�VU2&�n4��@"~��?'?�4�G��s�S�ܟ��>�&-�;Mb�K3:�|�����<>@�[zF�����o�/7W����h��Qܺ<��<�IF��P�����y�L�?��~GG���O�A�蝏� c��������K�r���?���<.@ī�σ��w�~���5�Z�����;��f�?l�Xs����gS�x�t��d��ˆ�4��;�$�(�E���$��ǜEV��OȡwH�4"Q�1���'t�R����2�����J������0$�˿u,F� ���69��A)��7o���$b+�^���5#�GM��C���=O�C�Y��2����s|�>�������`���U
}����&�Ǣ.
n�H�	���h!�
�
SG�/$X.�':c�H�.%ABA������b��0J�d5�IA4iN��>��*��N��i�h�{yS���2�B�%h��݅�)�z{��uΑ߮2DN� 5�ϣCp�#���f��rL�dl�%p��೏x]�D�hi�#b�9�3���yP��XQ�ZC<�K%����ᯕ�0�)q�����W�����t���f3߅�?dp�)y��[�s��|�<w�&|_�h�ux'�:[1�6w,�Z�����|a�)c�������Q}��^�+�-��?���͵E^�*9WXTԘ�Wa��zAN!�a�Ԋ1�瀱zR�1s-YLR���t�ix����������\Bs�T�D5��o17�f	MS�ޥ��`U>�G��3t��&��s柍~u�P�bc�M�ּNgFs�V@sy�]ש����`I<n����s&!)͚P%���dC�<��s����8H�D�EG�*%	h�A�Ɋ6s�V��a�\08�W ��>҈',p�9$耆I�A�L���3��;��a�7'=��	��c�u7��� X�4 �0;��i$O^�wh���6�$�?��?Q�跔�2r&gOT�L ��@�`s�:�I����k�
)��������p�ha�t_K� +�Q��<��m��(P=�`�b��7�Jg�#:�_�]:�gt�1-a4�P�_S��Ǟ�Ha����g��t'�C�m W�:�U�&�+G�b���D���Ë���|����ñ?��S�����7��
s<��"��g�؀���.%g�O��8Y߲_Ju	�,$��"ܾc^�W���&!ld̩rE"+���������i:�htoa�-�d�}(�o#)3�G`M4yn�/�>���8%E����4[��g� �b��`���L�UJ�[�4SQ����d8e�0~3gP�� �F��ŷ�i�5�Ov�o�R�����!�r/Sү�1>��_0��,�P���t�E�f�0]°�X"�W!ʬ�rC��㘍r<�Ew4��J���d�
pѽ�|�Ö����3PfUT�,�W� �풭AG4�u�>(�J�&��Ҭ��t{)T�UC��y�=4�{^�� �'aF�S�m�fy�k��{O��m`^�3�7򉘀^������Ù��|}�p^��?L��y��N�6S�0)�F�6#/�ymi��4�U�8��23��5bV?]B"�����8s����� �Y���D˿e��$f�Kf�=��3r���Ԑ>'������G^8&]�t��/�,yD��?Β��r�U?e��C�m�Q��j<*<zM�ݟLH�K����af���Ib��l�Iw�w��,��T5,�o�R��g~��$)�?,�WKB��"OB�^3ڇ{K=�l��Bfn�j��\Ѵ}�ib`�Z�O���hs:�I�VO_C�����
	V�_W�v3I��7l����)"`�
���.���O��3ף��]�������$�K��))��&͂$K��� ��#����j_6����:��tA�V�9M���KD~�1���>��;����G�\�F�!�1�J��S/!F_�7��f*xy���_�`�'��r���>h-��|ș�0��]��[�塲���0�}̩,B8j����f�����V�\�e_���hǬ��9BU�O��XHgX-`�k����.�	9���0]�ߖ1������UF�v+_�F�b�_ߨ�%隣�Y'��2����흾\��X��pPw�X�H!O��mOY{��S(������G��ȍ3���.h��%{_�Y�w�5�5X��\�6W�ݩj��X]uJtg/�L��d	AdbyP�#�o�A��CO,��+O�Q��d%�e&*?ف�ºt�,���d:�l�3 �D3s.m���w��^J�q�̥�6nw��W��Ud�����xu�\]��V�>��Jc�o�z!`�*_3OleI�̏5WRN�^����g{�M�z�$�t�eˆA��"�nU
L��VYh��O=�)[����]��ォ�U�=�o�=�����x2"�NH۱�aT|rN��)�繓��J�.�9��}î����[���X2����\O���$3�*X�>x�i�;2��I�� �rF1�;o��;Uif���:���T�=iˠ��.�Ln)jZ�z���>Oѡ�j��1=*���6��]sj�O@��F����NzR����di�-���OC[o��J�5������v�ӏ��Z��,`���L���fO}f����=�#X,W������
[���˛�U��9 �y�W��+	�>�­���RZ�Fp%:�O~����.A�� ��=�DT��!�8L»E���P��_m�{�0�=���W�Y����\k�@����z��|if�ݹK�z���u>3l�g*#P�9��÷i�\e|G�f}J-r�^w�]��}����x����E����2�4)(�L��]n�L��C�Q�\c`(ku�q}��=���5��h3{@>�4��Mˈ�0nx�p��������gqC�*J�Ռ����������n��&XH�u��Z��ʰQ��(?p�܌�����c/�Ǩ�;��fm���aGR!���=EA9b��N���C�'qtK������$�v�H���9�p%����Ċj9�|R�3�|�8]�a�j�7�%e�,x������Y��I,�%�ib�Ri8]��Ҙ�W�!MY��:e�="�h�A��E�6ekg$����OK��W���*|�M�����|��n�,L��(d=6}��*���p%�<I��Z7R{�B�����u�c�e�1�$���"-[�ѝOvt�)����T���İ��'��>���0/�k|l���N!ʀe��d�#�o��m����8�~!w��/�$yg_�,	�VMV��'4���
��u���#�<��<9Q|޻v��Y=kF3����=�~���i�;.��.��rF�=����P��67���5����ȷ���3�m�CN�1KOp��m�M@��]���,p�l�A>�x���<Z-�)�-͞�<$x�9M0e��h�E|��Zh7���'1?����E��MaCS_d?�/~u�/�7�y|�;�W������1���}�>�w�CU߬�}
��ޮ��e��k���j~Uu��W��9#x�e���H��>ɺ>KY��B)�Y&�1�#��X��є2ذ������X�R}oY�w�̀�����{G�ZZO�:���K�(��Zkh���(>�7�ZL֬�;r��.�n���6]a�n����V�����VB �4��0 ��~x'�;�
I(�(�N��&��2��<S�a�eW�KJq_�L��D���_�(�7쇪}�I!���<*������gh|�ī��SH�z�tdwGU�$�B�y6�����.'��ڹ��"�����}�E�{w\SC���H+�ga�[�a�_�߇IM�m��@�����B��x�{}[�߄��F��0���,��#Ƞǯ����?W,�h�Ɓ��t*�s��S=�j�pޙWu��#����O!׬��9�)��\���Hf�c��6��iR Fs���{�M,Y����������`���9rȆ�Wd�Z��_#X�V�b���UE���J��b����U^i�*��.��ݰ\���9���݇�k"|�!;��P���g}�A��]������!�~u�p&�&��a��	CQ;�|�@mQ��8���"�+b�W�^�n�Ns6p�S�,g����y���iʱG%`��4Ʌ��,fv�B�2{��૛h;�)�#�w�K�ݺ���ݶ�m��s[�Q�g�"O�G4^���$	�F�O54��O�~~o�M:��<�}t��2p[uY�2$oPb�F� ��������"B�R��L���s;a�bۣ��@�c��x>�d@��GK���d/hh������*n��-5Ax������K�пVaBgb�MJ������#�F"ł(����3E��
����ML�an�m���/��4#3���<��*��:nx�n ;o��{�s� �t�@a�IS�By��ݾ"R���;�Q�w�1�J� ��vް�p�6ۓ��=96ӊ�ҊlC&β@����]����%����Z��>J��}�
V}��y�1_Nj��EMa�ǋ#n{е|O�"���!2W+�C�`{�)dQ��<J�d��Dvwy���u��ڮg���@돳�`]�@�����~���x�#Z-��6]t���ÿ����� /��� �|����7��8�٫�}|�<�j�񢀉q���js�"�v�G�V5�u�s�xeS�BD.
��7�P�E���0�0��0��<_&k~��H�Q|eW�Z�%r�m��=g������|������vgKnwln����o��s�ѹ;���jK	(��R�l)�����O�g�ddق�?*�S�����]E)��;�S7*c�t3�@�]�2�ʝ�����W7J���@f��`8��!�n��D�Q���.��To�0����S��v����w�eET�5���E�F��3�I>��IB�`'r!K
��4�$�}h��9�|���[�^���Yn d�K���0������$��A�,���)��t\_wuo�Yl-�9�G��s�w�T!�M?u�hJը���9��C�a��ǵXj����ת��j�+����X����8HL.���s�b�C}(�Ϭm셉z>�,Gg񫣾m(�g���bYGG���3�}x��Ëo^��Ë_�ˋ���̷9��8��ߚK)E�/|DE9���%WD���uoߟ��ߟ�������>?������Ͻ}~���so�������;A�>?W˧�}~�;���FeR��
�m\Z�r��<��xeU�|%�o�֘�:~������>���y����Z���q�'����	��"ķ��J�W׀�� ���M