XlxV37EB    1dd1     7e2xڽYmo�8�ί���
]����ݕ(��"u��BW�N��$�v�vh9ݏ�;������C	�����g�Z��*�j���O�Zx쯘���4��I��$�F�ǋF�� ��ۭV���d"����R���t�#R��Fz�p� T�*��M�X�M&�ǻ<B�2Z(>��r���@Fr�C.���/�:�!�34QL35gA���Q��p�51��_
C��$R2R��U|:��hxc�f�p)��wZ%�V��Q| ��b0EB�3�+9�aVm0gtAF�Ě�=x��8�VR�3~(��H.H+Sa���L�fz7쑒9y�t�Nc3��<r3�S�w�ǎɀ�q�Z��g�@�0��B�#��(�0�d*	��n��·��Sc�4DGB}_���I�^@�S��.����|��:�})�A}9����I�Q*��x�B>I�'�Uf%E�W�JtER����G��'i�s���O���)��`eɅ��?��
���,��䑧�4������:f���n�H�K!5N'��rMx�(f����)��3��Z�� Fʈn����\A��ఄB�T;�1R��l�c)i�$)y�"�4dJ�協I��՗��lG�1nçQ�ЏP�R��[��Z�Ӈ��.wW�RHG!ۆgK����P�0l��_�8D���#?=4-�i� �Pa�,a���q��G��V���Z�Ie����s�;f���G2Ag��z�g�������x��s����/|�$W$Ɏs��ٯ?����bی��<������f*U{��mMq�+�s�d����kO-����˧�IQ�{�D���T��ۮk���M��k���|�
��ͥ��������J1�>*R{ 
�=�P>�'P�u�0CN�=q������s�����?�L�/��W�������)6��S ���~�S��e���y��I��ؖ�����n{K8�)
/P���]���j��Ja�i
v~�Η�� %�ѷ�vr�1�x�B�?h����Ch��0`��-��/&'�0�벀���ct�e��v�c	��(6�;�Z-�$��"�W���+���0��.�9�"��9�ӻ(bʇ�(��$6l"�q��K�7�CI�2�]@!��0����o{7����{��޾����M���KE�G
�	I���]� ?�]]����^��ӛ:��˩�����y�7^��Qg���n]�GC�6Tb�=����eV�r	����������M܍����`S�2���j[=M@��w����������
�O"y����Y �+Vp��ӹ��1��{��:`��l��֬8ԫg��Ĳ�[�q�}���F�	�E����k�o�ۃڵ͈ASA�Ι���ϗ"Oc��m��?�b��	 \q�h�"j�e$�u�rѪ@�:�Ky�%X��:[M��3�&fz�Z_��X��R���v���Wҿ�g�y��z���m̉z5���j`ˌ5�n�;ݞwM�YJ��3���WR5�����eVK�z	H��=�FV�+�E�u����J3���w����KӦMB:b��u�����'u�r�6�^�ڗ �9�bU�N��:�bK�&����b��z��1�<�� 9�I���+�w��p�Y[W��L�}G�_�5�q�<Kjq'W�q�]-)�a\m`\�Xm<t���V�]��)����y](�T�b������/uA�(��il�q�h�u%�������O���F��y�U�_\�y�'�^���)�]R�7D����n��ܢl+Ȓ5����6��N�u�O�we�+��7 'Wf��s��WK��V�/��DI˂ׇ��c㬺�	���s]��Xt-��GLݨ�\,�n�Ճ<(�!�++��/'��"�\/��$ɱT�ٴ�dn��,�d�r/�Y*r�#�Q鼭��:��ʴ/٤r����~+�����A&�`{��I�ת�L�u�2���0�,�_}s�