XlxV37EB    1c99     6b5x��X[o�H~�W�>@�&M+AS�'k���n����	���h���gf|C���� ���Μ�7Ǵۖ9����_��M�}�����pb���v�)�?�_���]M��Q�?v��u{��=�3D�D	9�K�p���Ia��m�>g��#	�Ʃ�W!=�������O ���-d���c�kL��@5`�y �4�ᚺ��L:FV��G}���Ć�#D��0b��J�Z�h�����%O�E�!ͳ̙#׷�}�,�d9���Z��1L��Kfa�y_���"�o=e�\ѝz[;owτ�5#���H��Bdi�kя��҈��5�����}�E=�����~=E9^���P(��Qo��e���䵞%M4�e)� Ж?�>���U��}����]���̧.�%��|�to�ȥ� ��|���RoK̢J��
CL�(�<�	3�,%F���`�.ْzҿ �0ϱ��y+�A�{R8p��}9��:>?-���̣���P�;���P֪ x�`ŗ+� ��e��t��N��S�(�ɇu���Ρ�0r>�d��K:$�9ma��(��4�����aY��._�z�	v'QZ5�Ss�d3�'�^?���N����B��]�q���ptx�L�0�5q�x�Dܵ�e���O�y�T��9a0��?�^�5�&
��ޑK�ri*�B)j�����@	g&>�,bu�z�%��{�@.u<��:���$)3�MB�[~����Ƙ��ڎG6�$��}򌗞�����o��L����M�����(�U=v����$�%3l+�B���9H�1��_(LFwCXb�N���̃���?􃺘���A̰Z�d|Y�����{��(a�������]F�\F�q1b�#������K-�*3h[Y�|��+�Fk����O��N�SkSID=|yH�XZ��[V�%�`i�"5@�g� ��=m�[�^���	.�!�h��hjF���&��ed�9=��[S�O�^�XT���4j���z�����I�/�Z�^{q9��]@}�D6�y�îlӗ̊m�]c����auÙ�T�ZԳG��N�D�ʾ[q��]�81
c�Be�������,V����~���_�����VY�c*g+�-g��-FY�5��㛾�φ����L�rc��&�96E���#-�ᱮi�X NO� �6��O�i�d�;z�N��#�	.�Я��$�{��*�:^����p�><^�'�8�c�F��cZ�Oڴ�A����)��6{��'o��=���1��K9V�����{�;J�IRM�>�M�z!Y-]���1��������L�Q
|Q��L�z�o�m�k�N+ث�R���w��|n�*!�Vޤ�v������2���Q�M��=�Zo(�Ŷ-ޮ�������[z��j��wR�S#�6�����	�xs�C���$���!�Y�k.�{vB��A��-��#�1#4�M�'�L<5�؇�v��۷$�Ed��"�RY�l�!�`����jHf��f͖"��>��ߐ��3����JզfiO�}� ˤ0����>���f-��G�C���?�U��������M Ҹ����9y=/������j��V��=q����q���%kH���KU��*[e�̵ۜצ����F�-n�c��w�x:2&�G:���Py��:��p,J