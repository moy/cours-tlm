XlxV37EB    6f19     f07x��]�s�6���霥DvDIv\��MK��~�$����á%��"U��s�- > �ć�kRi�H"�`����b���ë}m0�&����@�a8;A�--�;x|���t�#�ۇo�Go�jK'�ݓC	���������\�\h7�������[ݙ>�zKo�E�h��:�!�{����d����BCkz��d�DT�Ev��g��J�61�Ė>�'Ax/!~Ŏk�VX���v['E�؝:������0�.�Q������Ntz��4��:�M�k�9K�N'���� 7�y�=�Nd6to;�EJ>�g;/'�W�2"�(���CRw`8��~C���u.m=�(�-�$��>��G�L�	�ƽ���	J{�֬�Pjj��/�Ljj~�m�7mf<�
>�zލ����WDX�(�7�K$�-��<Q&�h�9�%)��;��3�,p��'��>'	y��h�C&�0���.����͔�.�#E䦼�Ԟ���d�f����=���t|�f�w�c6�A�^	.-Rs՜쾞Z��[@��5q�0�(��3HkP=�8@����b顅�'gD���1�0H+�A
��f�+�^4r��n�rz2�t�X`g������S�x�F�:�V��8��"n ��t�N�h\����d8���<�~z���͕���SŎi�:���~�t�~:p��f���T���ށn�\�����Ӡ+	�\SǾ5�?�����mMgb�����4!��4���~?��3]�5�35��.l�k̙V���1�h�kg�V%�:�SSw�4��������5v��(�-G��8'�}�����3Me�~��q_��otA5������=�����D�����D+���K�=F�ȳ�Q�T�vh�&����w��ꄶH2�����E�+��m�+��=�V��E���B�Ю=ִ�F���þ�D;UEI��� y@�U!��:ؚ��x�o�9��\xgc��z4�TI����V�P��fnc>��z���h@:�#D�IƼK﨟��o�TV�k�?*XyV@sT��i�8b�"���uazwX4�T���I{�uc�nq��<�Ѝ�SM. ��P#LM�\k"��!$���Q���"�40�[1P�Қ�`���[�/�2_���	�$ax���@�] ���C��8���R�m�&��F�l}�k/�D� �����*�Ʃ:Z�
���vv�i�%��r��gJ~��iR���D%�)�uMSͥMj�l_:̕�iӗ��D5��uO��,��?4�>R/�W����L�:�9ЉH�CJШ|��L6���Fz�+�#�
����3���I�;P�	��r��(��3�@���YX����+IG��� Z�@�B:	��I�^�_�NO�N�I���d`����T`;�k71��a���Y����H�2Q� �'ؔ���N�k@�!V;����}���m�K�ߚ6�M2���~��6lP����h��ڃ���bAl�%��X�lv��5�/0�6����5F0�f���hJq*:e���
��TȹS!gNEu�wD�w˚��׌�Z$(�"A�o����#S�Lpx`��i/\����:5 .��Hv98�4��5 uR C�M��d��.� � ��9�b�#�T1�
� 41��������`�D�n1W��TM:x �q�YN�D�ճ=�n
��Ki����a������"3��И��A6W��X�\\����~&B+%�n��|1`:��M*���ⵞ)iZE�A\��4p�0PC[��%ҥ ���yg;hH�u�1&Ĵ텐�%������jQ�hcؤ���ީP%�g�2����A�fL<�M�2�S�,�g���(l5��g'����㑑�ff�*��(�~'�5�5]-�t	�K�L8 \ߐ󉳲����A[Αn��c�ʓ��� Y�7��`�g$�=�-e�������,w����Y8n�G��dlA�lH\" �\�i�B�B��4��"�E��������َ6�2F��_�G���N�ܓK����EcUM�n� cƱ3#׋Qy[6-�>���	0�8�ɡ�<ǲ_������篤���DXuʧ�S�v�7��Y:kC	,}#��Й�����D 0�L+��'������'��n�Ω;��nץN����#}� �D�T��B�EG�U��T����ESo5A`r�O�v�ubrv���N+���W#�����	j!l���j�[_�e��4�L[����䥲ɨl*�v~OU.oT��hT��Q)R)gT=ōz�]x��Ҩ[�wK�n	�o���ʤXc�����Bx��Dj�D�_�2G��V�	�8��]Х�%�R��ѥ
�lk�ЈE�_"�u �J���2m�;M:e��IҚ���R�1b�i=�HxC�LA�+�|�O��S�$9�$	�jI i����e��&����D�ɸ\��Ie	��UDƖPX� �
��gz�z�0��P�J)pj��R�R
wJ!2�>�r���Q���S���ޱgu�`>�����<��~_����~�8���{&n�l,s��C�����W�`c�+��K�{�:z�H��?���v����޻�w(`��U�H(�_t/�j���+�jh��c���fq���N1b0���gR�}B&'X��[բw��I޹&�:�W;��3�~�pF[0��8��5��&�<W�͇�o��LL�P����Q�VI9�M���%���s/�R/��Q�hK�g���D*�{�ݕ?{�$�Ď-�h���z�&��Q�M�R.��"@Z��Ti�[F������h�������B�]��Ǽ��F`�D��p����3�:j�ߠ�d%��]�]ڃVS�W�Tw����y!G��z��Eԗ����?w^C��':#����K�;�g�:�)�z�.�cT�uoE�$�c���֤z��
pU)�`z)�����a�C0)�az)�U���k�m>�g�$����'D��C���b2V{�.=빤�&z���h�H(!�oA�g����H�uH(Dդ�j\܄����9��de�8�b�ޥ�؇�l���9xxFb�>�����v+�f�Gf{vmx��L"���ᨯLvÛD��9�*)�h�yx勖�/�\Q�*ݻ�������y߷cI>I�c�E�!���qg�;�{u}�߅�4��#^�;d�'t)��|�(����� jg�O�M\� ޷Ū
y��\�<@����.��
�Z%c$ZI�b��י,j�J��?y��Zϙf��U�1�R����@]/K]�;�T�Du"����,F�U9�̩;���`�Pé5�)B��-�.k.��᫃����/-�g�ÔC� �[�Nsg��/s�S�+z�?�!�ԑ�WElwsV����j�/k�W�.{�/{�K	Oc8�e{�N���Y+�F��+B {VCV�#�{n%Y����^F}�H�V1Y��xC�B.0��	DEd����R�Ǌ|ާ	u�,��2YJ�di/��*W#����eg��R��̄�q쾅�[����塢ȟ���E�hXn���x��e�b9ٚx�[/V  K��2ذ$,����� �I(Հ�e�_*�ΫJv[h���*�K�r0�L+q�5q�Բ0%�v��v�W���C|�0_=�W��C~��_=�W�UC��ԕ�"���
�| X���``= X
����`."����cl��|ğ����'��O��$~f��ϢIOw�~��cO��6����ZO�OԅU���@��J<����x0X�\�9����0�Ib�a?(��%$&>?(�l���A���+Dtx����+�3