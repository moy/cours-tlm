XlxV37EB    2782     85bx��Y[o9~�WXt�B�jwh*QJґ(��TIW�eC�3�g�I�?~�=7ϕ4��H�C��}�}��g�lN���h�/�3�_V����>�����7���5������Cک�ڭV�L���m�j����^!�#�K�����16�	���ɽ�&��Ǽ�3��{&^m9EGXU,����|
���<r����-����@�m��b��e!)�"N]�wtq*G���c��Y�&k��{H%���r�9v4��V���w�59�x�pZ�D�i�-g�L��wG.[��B̕���6N=�����$W�18��?������~��l�<���#�����{�Nl1���G�H�ɚ�+Hx{'�Ա]=�1���r�u�\�UO�]��L�1���R���ڐ_x�v/���8x����(�'��%�_Q�rf����|��m��т.�M�{��b�gw�CE:�Gњ@��)����s|�ʙ[�!9� g�r���3�@�0��bG	9g�n؆Z�>(XNW�f�f�<&Ԁ��Eb��-f�I�Ĵ��tZ@�[�LXl�*�1���&;�;!g�����zh� �)r,^mAw̤`�]z��9�[@��l]BTu�<g��̻G7��&q���;&u]�O#l�zr5N���n[�X��N�hZ��p<3fw���_����f<xs�VQ�؜����pث@�ȧӸ�kګ�)��^<�3�3��7�w]�ja�Kfߟ�Wo嫙��@�b��jMЃ�Ę{v��h���l���}�|A�r�z-�pAM�p?B���O�$��!������Z%��)�F��'_�����Ƨ!���-�jtYQ�E��^u�~�:�^0}֟\g�YG�3��0Fw�ׅ�E�zn��Wz\��I}`٪�e��%�m9V�e�G�J����*�)r`BWxF�l�X��Ҙ��rf�q���-�PwkE�&5+ =�����V��V�f�+M� /P6н��l_��.|C�>m���p-�w*��K�B<ț���O�0�z����j�
��� �Wd���ut3���$;oP<�����!��3/$�����V�ϑ���Q~#W���խ�����vz0܂H��u�6w�g��ju��d�t�K�W!�g~�Pzu��� =�pd��FFWi��M&wl�W��e��`���UT�/&V��8�V� ���M|�%�	��O�Cꗚ�{a��p���TJ��ƅ�/�/�"������9��Fu�V�X �I��e>v8~�V�@�S���1�o�uA�s���M7����tS{��U4��<6޾���7�"�X�<놕�" d�9�'C3�2x��CSC�ݪg�˛���>�{��'j���%��WK�< �?�'.�td�9��-��j�Y�D�R	�uI=,�8��f���0~�&∍J�=w�̌4�E��P ����H�mV��SuA��#P|��4��v$&��& `G/[/WI�'@�":�E�g�N���"��x�(��_k�kҫ&��s%8����y�9K��'e'�q4E�%J�'\�T�'N	:ZB�1~JR���T��-'B��W)�}9*�~ۑT����,�
{~��H���F�X��+M譇���Q��U�~g��~�/:-�]�g��u}��D�U��f�ʱ �ё��z��4N�k��;�xe��T�x{�zM��{aū��%g�^;��P�<6���IA��:[|��K+V�x%#�td��V.ۿ�͵��������F��TU�i)e����vR�H��+뤔��-U���CQ3MCdH�0��C�{�.��~���#:-I�=�I�4~��偤?"q!8�@-��6�A�?pA/I��a���`�q�>��f�c�/��ý-%q&��Of��adO�����@�E?��g�=ǀ2�����O�A9�J0(�)cQ�(a����H�G�R�L;��M�
5ę>�jM�&���*t�B��BgY��6�ڕjk/fC�{�uA��C��c�W��l���Q0(�<0T!/�AM��h�?���I��Mf��f/Ⴆ L�ß|��l��x#���qk��R�\2Ej_ʟ��;�\E���]��%e��j´���s�h��������,j��	�|�	1���_A@�������h韜 �����