XlxV37EB    4730     e14x��ko�6�{~�-n�='���p��[��ĵ�]/��Ȍ�F�Iv��~�͐z�)�i��5�8g���E��x<��xٳ��5i<8~��#�f-.i�3;�>u��KN���暘'����������-�h�?߉�9�=-�w�X�5_���/!Ǆ��<��^OW���8{���A �p�y���L=���d�'D���}�bјFk:;a#/Y�>���|8��֠��L�������pp�Kc7�I>|P�$��N�,VOJ����8�V̦Z|yF-��XJ{�܇Q!;2ar�ŋ�0zn������yl����Eq��O�r^0ָ'� n�s��[S⇏$����-��4��A#�r��}�G�X���h�/{��d�yjJ�ݓlC$���R��i@#ϭC�������=Kf���$�K��|�u�0��I(Y�c��Ч�?j)dk��U�:���xn���L�s�A!^��ޒ���01��Ͼ�,���i�U���t�x�ɻ�Y�ӹ�i2.�
�y8 �5�̷���*!�0JD<��mFמK�ɠ^��0�X��Fk��94&� ��<z�=�Y�gq��
ԢХqL7Q�eGם�x,�vh�E���t�-#�ػ�&_���o�ۿ��������n#'z&�^�w~ ��u'3��k�懳���s�O�����'��g�a�G�>?a�.أ	n7N���&�bo����)�\��jF]ȋ��__�<��R#��F6�F^|�{-rx�L"��'�}{؁r��7�,�E�C���4���|�y
��ju-��氙���N���ǥ5 h�DS8h#\B��(��pz�No8\_��nwd_&'�#�yk�̀W��ht3�lܛN�ѯ(���	;��o�Ч��\�������v�}q������Kod�Ҿ��uU�!A��q����)�bݜ�EB6���g9W��/����M��$���Mm ������ѣ�L�Ce�H�>�����H9�ω�z	{�djR��G�Ñ�u��u�3KE`Q�,:|�͵�������Voe� ���y�v�ɥ,��0@F�e����PN�S�ÈiLq!�V�c�U3dw�C�v �8#Z���ߎ�:
7���+;}G�e�i���:�,����
r�����4w�L-Erpy3�x���%`�W�]���@=�=ӆ�HǏ�>���(��:#fy�QFM��<װ�`l�Ĥ'&H��U�Owd�p��X���^�;��lWy���GN���Y��ζ�է�i�}&,��p6&������԰��5o�n/���2r��'�}�$����D�I�%��uo*"�Mk6��:=�H�la�s� Q"��)$��0��0�G�]:�U2�vj{J6��5��n`bA$t��̼���~�I���*`��1���&9�8ќ%��2�Dg���LG�����1��r�?�σѤ7����Qy
��I�ip����d&7D
u�<�����.3���\Z߄˳��a{4i_��:�V���k��^�G#�q&am�4��~A�/�Hp��Z�ꞹ�|Z7�ej������ ���|�C�D>{QB�,Y��}�֡8��'�{c,��/Ɇ@/#���	?�C����ٜ���u�fN�hH ��G6�ݻ\�?������U���ߨ�݉L"S ����k��	?
��P�rd1�� �&YM#!Gr�SBc��iZ=Y6�M}��,�F��P�ӣ�R��Ұ�Ѡt�����h�B��i�,;K%,�~6+�M����%�3�բ���O�U��TR�PȃR�D�g؃:��sQ�ːPXG ��7�~��"ۀY5`aֳb3nG)��<��X5Y?IEP�3Ӗ��J�PӍ�H[��y��f���`��b�)������E�$����Ok�_Qr�e�3�E4�Ye����F��]�3ua'A�?N �A�o���P��Wy�ggi�I�ɵy��.�������y�1)��_�����R6;Bc��i��)���8�!��E�a�i�?+C�i�{2�Yb�:X���C)��p*���0��/Q�����j�YwS�t�ަ�7ݬ��f�Mw����L�b���[Ѕ2���4՗C͏?���[.:~��~����Ҥ�.bS2�nKsK�aIR�VU�(��
�
�,�V0���P*��V:����<��H��Vr jv@$�USE��ё8�~�mz�R�=����+�}t�s�X��b�!vW��YJVp;�T'Yw����x�4Ikj��p��^t�!?�m����������fx��M{t��G)�3n�k���G\(N&5�%Us?�ι�����sw�Ae�GM��0I�� 8@�:Rʧ���*�u	ޣ��d�/����׵F 9�&�4w�%u�01�e�tȜ��L$����>�5�u�iw�=���;W�w����OͲ�W4_�7��I�^�e-o��*YEs�)���ݞ/�N�^��?�R;>.�M�����".Ï� 曵��
�;��ĔI���w{jc���U([E�X�VV��7��v��R�4�S1)zv����I�F�]��N�{eroIKzs�:mU��,�{ʼ��@H���[rF���cHf��ew��FELft	���A�5b߂yJX5��9�P�����a��wVĦ~Z5�� V��Z��Z;Y!��cU����ғG������C0��:�Vj��:y�E�����F.%N��i�#��|~u� \���ʥӎ���4��ﴉBa�͜�*[�D����S4�1	1�� �!�~���@p�P��cBn��73���ӆ�rA��G��_���ȋ�̪���"d�y/��m®(��aῐ&��ӮE6�	��W���ȯzԍz�a��Ŷ�)��V����*�������S:#�*K*�ζK��vI�,��פH�Fjn�"�u�$��[�H咾�0��j�J1�m�|������6����`#��00q���X	���C���!���H����&��;��Ɛ`\�T��>҈�;��c�ȡ�������ȯn�Z�;�i���c�E�����o}!����v����0�*B��qz���4u����N��m���RŬ>�,�_��p�J�6V_�h*_�8�����B�m�Q�7y���l�7����v7f��*7l�<�,��F�ڴ���x��(����j��aR�S���������`��/F�L �*i�E=$�����޳��<�#%�}ưoY�3� ����x�uK����;){ �^������N̾^��D	Vw�Yn�=���
WZ�&;�Xyf癣mn�����j�g3;���Y�"m��"�""��3*���b��Yo7���F���~��s�-����IS4	���2+�.im�	�v��bTM'4=�ܮjm�	���╞�.MB���j�cT���A�J�����]\�Catzٻ݂@�~�o$Jg�Lr�.�$�l�9J�lM�GD�4�A�1�8�L!O�0������"�