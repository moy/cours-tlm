XlxV37EB    1cdf     69fxڵXmo�8�ίѕ�"�	mW'�]��A�o*�DuZE!�`mH��Pz�c;/NH��"�Z"�<��3�̘fs4����[�!��nj��>8|�:���[�?��5���^�k0[&����4��m0ڝ������C�M ��0j$��|��@<N���:ʉ�W!�
V�o=g;�\��{H��RoӀ�素��s]�!a$\�YK���IU�d@]��K҉m(������^���2[�I�Ҁ'��e��%�����Y�� jr��Kd�)Tz<\����Z��*�����S��ڞ��2��e���Nͦq�4�v@C�cOTdཽ���[q��$�e;��	���{��:P���,����w~�&(����7�5����hSO=&D�?2��� ?Ж�?'	������֙F[�taF^�Gf��R����c_cbV��6&8��G6\}�)83V�sVa��(�"��y���R��P�����_jĀĕ��C<�9��ܳk�g�A��(����}>��9?ˇ枩Kv���D[���k��Z�V��ƣ�j3���Mz�]�,��ǂs�|�r�)��o�/�9H�،h���C#�fD3����Qֵ�S��Q��h���?�_�oC�������oO5�NC;|�a����P ���,J�����e�n7��Q'����/�֗�aX�"nߒ_}�_����D��et���=BT�EX͈�ڡ:���ꃶ$�jIʂ��p�5v�O7�1t@�X�����E�nyQ�Бb��8����7� ��ኈc<�!����)��ճ.I��+��~�,�Y.��nj��C�4�$��A?��s k����}0O���9��.R�#S���]b{
�q��¤O�y�p�V
́���AqU#��޲3�T-Ɂu���E�/	���14�+��Sc��G5?�U�+���y�<�T�J��B���q�{ݓ��O=�Da�E6�m��pB�8@p�,i��\�G�5����uKNOOw�R ����i!��;�����*>�̖gc#(�>���Icv�L����a�S��W���ѐ���5|�E��T���ۇkK��f���-9$Z���αg��-����9�˯�'}"]��0Ҝ�>;$��m�D<�<�Q�@מW����}���rӕQң,Y(J;��׽^���2B�29�4�n���U=��L��`QUD2�@ꂛ���V��aTE	�.[e=�|�뫆\H1_L*J�Q]N*�j��� #��荰�`�������yP43�M�in1=�'��m|x�͐y���1�i���x|�j�@�,4��L,�)�,��p�'-0@��=�F*3�	�\UZ	'"S�Vz�5Wo7�ZdZL����.#�����j�o�\F����i�F�����$��H˸䘿�iN\'������͹(�䕟bǕr�Q�̹�k��Q�4U�ێ� ��rB�]n餍�^"4���w��S_$�2��G�Y�Y�l�X�9�Fh�@�b9$�V�ND�B�z��eE������� #7!�"��j|��#�RH�_�������F���/~�]��ɪ%�������u;_�±yo�&s}'.#pl˞k�;����0Q^�&y����Y�Hbf'�x���2�O�����G�Lt��'�|Oխ�.߰