XlxV37EB    5587     983x��\[o�H~�W��Ji���4�hJZK�	H�hUY���F���j�����cc��f[�Ф>�9��rx8R.?��3��?7������E.���O\ufZD������8X!�HFX�:oe�-�H��w��1�|��4�G���c��':�'�h���7�����ߙ>���Kv�5�=��/� Щ�xr����&�eڏH��#T�[b �wE�#F��H�P
Յ�=�nx��Е_�뙎-D+�H�4J�D<�5~DVy �zHF�93�ߑ�9�̅"��G��d����w,��.N�_�w���W�)���q���x�1�~*J�C�]{f���aG��L{vn��k:�׍�龹"�r�#Ϝۚ�u����W�f��-G�/p�n�7��0W���_=6c�Q�0IQ�����&���A9�T�O���� 3�&�������A	Q�'�A��fd�G�?�
d�����:P��I��<LM[S25�DP�<$�sA,v?Ǎ�� ���b@�UjåMW��Is_����Y@�Z�LJ��t7X�V�hdq��b飅�+�3���2u���U(X��\k-�a�C<4����ߡ�ł���7�щ�u��ë��h�V�±��-|�S���\����AQ߿������ó���eN]�}B�`0�5�A�oG�o��37uU��;G�e�����:SK�����*I�Ɓ��G��G�hLݍ3�w��M�|�p�{�b!񚚕AtKs���_��
H��hDQ�5�~O�l~�Q�_Գ��r~�BO/Xr�m���e���tO���T\w��`GX��.M�uM�4}B�l2D��C����p���XyHc{b��q,��|��.ԇj�0�,uu���I�wP�ŗ�(e���r��r�Hx��D��,-�ட4_�]��tvv�ұ���@EF�/�'*x��O^�<��$��\\��_�5��:]���ΣJ�6�k4B�E��HF�a����O���r���f�D%�?���R	�/�q�]F�]�zg*!�eD\Fl�;E���*���R�ϫ�W`Ԃ�%�d��Pr�~���&�x�ǿ����x.�3�+�-����q;Tx��C�+�
Mǐ��tAs�)I�`A�7RvrUxK�P�J�����b�W(	%�Gdw�
�^�6<�:-��J"�5X���f�����*;�@������h��P���w�j�>y�`�fr��V���~	��)�<4 �D�l%`��B��Xs���+��Z�&�_-]hA�1�����+Ӑ9C1����pܿl�h��$|U����Ӣ�K�F���me�kby$M�4�ksj��4��"�Vai�ѧ��1hH����z��M��@L7�IA_1F*cZQ�	H$�=Z����Pl�?�qK$-�����P��n���P���*�j��oS��X��	��#�n�Ń�������g��tO���[y��,J��xB�>���@�*������Q�s�@���q�݆�$�`D��E��I�*o�xdo�xd�5��Y=��-mJ�w&��[�9 #yH�@�z����R}�^˯�w�����Zz�$u��,lį�X ܋T�����u�)�w��4^�Q]X��S^��Ӹ�ݓZ	����I:��q�����Iz'O�$�z�Y��ǋ�Yΐq��3�v��ΐ;ir�h�br�X'�1�#R+�t��҇���q��q��q��q��q�ҝ����9u�\�tN�e�dQ�,ȑ�\�u���D�Ai�Uϝ�L�_�Ŝߕ�3"o�<+�c<K��q�:~Ēu�"?\�/��Gm�;X֞���Z Q��e�~�����^����p�.%����.��^������W���Ϡ�N�m���y��%AY�"SY�F�M���0<�"qI�^,�ė� ��M��%\��",�$�.J,%.8D�5���IϕW�h�"7���J���:���хRt�|+q�J_��v� ��m%�'��&��'�%匧=��!S�A�{���[�oe��Mu[�okCZ�JPq�V	*n�*A�=^%	{zT���+C��*C��	*A�~1��$��a̷|O��pZ���e���g(����g^��$�q3����iD>��nK�]6�l�����6���&��~�%��x0������
n�H%��\Ɗ\"�5P�{u��qTK�x�F�`Ц�M�ު%n���g_8�d[(�\�XWI�P���G|�}���G|�e�go��&Q!��m�$\WI����>S�J�^h����O�x���O�x�^8 ��;�f�]4'������oW�zH�R�b��L��7����ݖ���z�ہ~I��Q�gu�����ճ�zVW��Y]=��}���zVW���Y]=��#~=w�gu���>S��~�Y]8��R������Ej