XlxV37EB    14ee     651xڽXko9�ί�J#R���Ֆ>���*R�V%�Z�*���v�gm	���{�=��B��· 3�����Zz�Z-��=J�������4mΩ���Q�s��}rtD���ӧ��3r^8'�����k��gӯ��j����NI�d��L|ae-.�Ç�J<���VM���o��t��o*S��I���M�QX��J'�\�mڼ*xrU�Χʑ�מ��P�QnMn���.�|w�R	�Dv<���΄WF�oz�$�*筺,�LY���
�JK�J�v����60�!�3��KI��i����
;�ꉱL&����lAya]!�'o�O%t�3w;|4�JW$��J9�dt��tS�;�}��^�I՘}v������@L
a����g�XLk��.�q��ܰ���'�3�HcS�'K�R���J�o�����1mnrD*Α})�	�Rn�%�fw<.35)�O9w�U*_#*�"ύ������{������|&7h!-�N�w���a�}r.��J��P�)Z��Z��҅���})>�	+������9����-xsi]��)"���~Z8x�*�&����c�F�4:MXi�m��Kцe,��Bh�i*�ӛ%�e�v��4�ܱr�n$B3���
�l��[�݆��������ËV(.3�/�t;��aQ0r�@���8n�Z�7�G���J.k"��Ҭ A�h%W�x\��]�ٯ�8�*.*�fҵ����~ż�NeR���-�W'�r�y+]bUΩ��n^|�+R�5,�����ǿ����"c�m�~v��	�)����zω���O�ȹr+�p���h�TE�����ms�~��(5c��n؏�A��u���S��5��/��L����=�9��
��a�旙+rj���z[+d�p��VV����n7�VI��t��j�h�����:x(���R�pY�O��V%��F���b�a���������ϧK�mJ�mYs�	�z[4s;��Z�!6�]R�K���&R�g��B���Us��,��Q��	�1��a����0}��a�y�]1�;L�?��hP|8�b�Dee?Ż�TP9�0�慧p0T��z�E��"�+ͭ���Te�ق+TF�K(��`z���&�*h��� �B��_>�O�����Fs�4b����i����|p�}�z0z���wg���*2ui�NH����5�G��v>ef��Q��줍�E�&���oc���*��5�<T�H���"k��E�˧=�*����ֻ�1/[��(��n���e�����6�s�9�'�\zTh��Y�)~o�Wһҥ�h��3ga�?p�9MNf��v��:�~|�xr�@E��e���%�*�Iw���s��`⧇'�k1k	�v�1��G��[�0�cT1�k���U�H�q�|Euó��W��sP��n�4,���
��m�
A�z�{���;<��<�#��r�a"�g�g��\�Lc�M��ɬ>��?���!nK����?�67Jß����GF�.ؔ?j�ƃ���%���A��{��уZ��FyА^Q��
� Biԙh�^ �5�� �м�����o�1>|����06*�G)G}�j C`����D�N�my�|��/j�&�3�