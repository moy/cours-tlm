XlxV37EB    7de4    12a2x���o۶���D: q��H�.i
8����lwk6�	��$Bɓ�4���x$%�Iɱ�e���Լ;��w�����/��-��O�7�m��C���C����zn�	�}���Qs�-j5�o��w��:l��0r��	"d=��U�Կ�>��1;ha/r��o�`r�Fx-\�s�ѹ�k�G�����k���G�;s��:�{�]�G��f�"�(�!�t��<��*f�ԝa�y��1y��_p���@���n���P����G�p��`1�/P�N1"�����Ѕ;	�����H�!�X�!RͿRȵ3�YD�~�uvr>��~r���R��w[�����Y�M�o:?A�G�~@��$u��9^FǑ��{���¿&��z��5c�;�=��)�9_��xF�-<�,�s�ō@M��N##������EH�r/lFT!������r��\���S"Xag*�O��<���=8O��U���� �u}���	���ǌ��w�3�����6��̟|6#0����f��������WO�(!(*C�X ?/)��p�NL��k��Ȭ�Zn�uLQ�u����n�-�ģ���bY~��W�
��Z��"�t(P	�Dě�c�s��t��AQ��0��Ϩ|ķ���q*3Y!�8}%=p�pN6_O��u�,��ϰ	�����'��?���/��"Bs��}�M�6ŏ.�s�ƌSO���B��Z����!�y�}|��q0q�CH���!.�Hظ\u��P�ڹ��� >�u��"��.G�э��o���ӏ��kw3w8�W�b��6���o�a4�g��;��ͷ{��l�t��̨�x��i(6�<�z�1xy�q�n4l����M�=�u�)����AO4鱃hf����#>zn�>0��w��F�6���`�S<�9�����U�9�n$�mo�u��8�ҕwGV��9<Fͣ��b��u��̶.;'�V�<��k�7�)�O��" �@�o��tF{���*��qhٗ֯�:����N�'���ϋ�G���54ľ�O;��96x:�6քQ{(�!�H�Q;��MH	O����i�?�cػ�?NC{��3�J�2�i@�2��;Yt���H�awNa�;q�)5��$=~�݀�G��f�(F>�R����2��w)��"<���#�@��#OόB���w�=�
��e_� � d�e�&� G��� "��z��[L�AĢ}[QcK`Q�f����h��Mw=�ɓ��T$�D�&�&"ժ�J.,/�)�&�FΝ�3&+��L ���'۟@Z9�'[��� �x�`17�h�({H�B2��1v$�L�2�U";B��l��p�QR,吥|9f>dn�E|��Kg
�ɝ{x� [���S��~�7�tw�'p|7 �c���QQ%č�_���d&x��g�g�ZMB�7��S�>!�'�*w�@l;	C���`d}jՀk��$e�\��^w��e[Cy�.��*f=?#���خ�A��SP���^��Ӑ)�*��˒p}O'��Q98JP'a�����x�S¥�b��W�8	�,�$�Yy�R@G�����]���gS�g��u��hbj�ի�NO!���Y��&z�w6�N���vk1)�t6�Ae�T�2[у�4��:.jw�"�5n�5�P0{21`��C=����@��z��`Ð#�D$�/"�e��t�D�H�_u�fl�?�P��7ĝ�io�vGRv����JRdu�G��d��T�^%n(
�I�"��b� D�do<�l�ͼ\�F0�d:	�	j��K��ؖYn����G{��|ǻݿ��݈[#O%�\i�o��7�#-�H��b@�b`xŴ_�b���⷗��7�o�e�e�Y�0��-�M%e�����:��Dq$@���=��'�pZ�H�o:*n�yNX�����=�F�m���a荹�@��0�ys^^�a>'<h�3��p�-r%�L�{����>�[�Hb��-�u�A��ƃM��P��X�e!)�G9��ݛ����_�C`%��1{�W��+j�ڑ����dpt��ۃl+N�m�K�������JE\�CY땒##e_���+fY��L�%��$�,��J�F!�ц�\E���U� �A�`�a���l��[��=�xiψv�-a����X���%�D	�T���4��ڽ�����mwg�k���a!�
6��e��[(�oa8�G�a(�31#�.m+�G��;̭��ns��5���v�[��|��Ɖ$}y:͔�ڽe�J�ߌ��?�����Y�έPpzs���Kr���jfgH|�@����g��b/�-p�y�GNpG���C�-�ͧ�;e%��O�NB�f;%I�.��n����ħ<�OZ<�-����?��֪Jh����^	�2\5Zh�l	�Օ��+!.*P��U5�vu�5h .��H��W�}�`��������p�W �Ƭ�����z���.�^i��P����Z=��U�m�jG���*��/��(��a�$�4v6�,����Ka>.ٞ,�l�K,��Yb�iM��{gG�;��b�*W"��s�;�Ñ=�M�|+RŻ�u�+��"lH���;� �c�k��(�<�����>=�ϬK��wa+�䠩�Ń�Z���-C^�1���*tM1ˡ��.}X��=�ӕ�u�ɿݚ�P7'��EU)�/)[k�=�r�P(y-�<8���O����ղ���i���_D�]
Ov�uud���$p�a��ˀ�(��0!� P��9�<��H�8;H�� �&v�A��|�Y3k��ͨ�L+��oh]f�ߤ�>�9��{���:��1�X��O�Fضh�Oe�=i����9��*�p�ٻ�����آ�ޣ�x��� Ӯ�~o��J1?q��"��f���!Ij&���:���LG��n�6<�]�q%,ӣ��5�,�ݙ}�	μ#
X��u��r�Ԗ:=����3�DD�b	�ie�1��Tb�w��"��7�M G�(��8Y)Áo�0��!�5����
be�T�(3����݀Aw�2��5��>��hN�ڼ��3�76zn'0���q�WL=�������n�l���9D��IF�QD�h�چ}H�:��Q����Ș�R�Jq��)�����d�o�VzȒ�>y�x�u������ͽ�-���/��^������w��?�6�E�KpyF��Q��l��a.}�]י�c��M��2r��	<��!3�$��}�]�+G���3�侾a�����bA>�q��WZ����l�TF�ܬ���7�i����0mU��
6��;;	��˫,��nk�3�\5T�
���UlE�������N#2ճ��J�Re�v8Pz_!�f+�U��T�hB���P�XiWys�{u}���H"z�|�`.����"}���7���s�Yee�Nk�L��ʂL�/j�+0��K�p* Z�H}�5�	���I�PξJ)C�+�H��Dϸi���RTP�ڮ�(��*���d%�.���O�V�eY��뷗[H��OY}�uW7�7�[I��3��oW���e�j ,�d��Ҩ�T5�vݬ�F�y�&ۦ�Z��Ek7Rg�̿l]�Ie���f��Vq(�R��M��ь�M+^j,/�L����p�d"�9�d���e-���W�9���78���H�� �C��灻hD� i�<����N����|g
����x;�/���<�{ʛI�RGE��?�L����,�W�F��Fb�p砇�;�zO�QPU�@�����B���-�.�Ȝ����\H�%��B��a^��>Wc}��ݛ:u"�2	�@��n5L�.�ox�o5�ƽ9FͤB)\iC��v�%�ǂڥN��W[J~��O����Ӗ�_�Q�ԗ����=~"��Wwz��󴭺 z��n��>���o7R�KZK�.�M���˥��+�{��-�� {}�IZ����rV(���4u��\s������-T��иAӴ#��<x�Y݋��ޒIWsf���]zQ��;��T�n�h��=������1XuU�k�0���.|���3�ĭ�&ni�֛�q�{����[�͊�W�=�m��UM
�i!>��'�Jg�;<ҽ�0�{���;��ԧ����z��P���w�w����e�,e%|������bd��%D��eϦ��#�*`Ɨ�.��/�L���:��
����gG�p������9|�q�׽V��kk�t���~��*LG�m�q���J�XՄWz��Ix��"t�X��υ���Ϭ,�����c��a�g�xA�҃���0�*z|L�*7��KF��å1���F��v'*F�j
�({��!Imi��M.�'K�
�?b&��5��8� y��^t�_ERx��)�#�[GEm0����E�U/{�ߛWp��(�>��sS�������<{w����x\Hy���B�#���|���3v���-s���(�ߎ�jl	]��23z9���<���l��p�Y�b����)[r{��zM���J�u9Iʿ�{OV��,|�5߭��	d1�6�l�p��~l�5��-;�Y��"���utl�!�Ա��;�[����vr�H-e[���VV�W!-Z��QW#L@I2Y�.kz��K>�gKh�\�Rk�3�+�7��[I��'���?���z
���F�v�\��Kr�`��${�hV��̳*o���Ya�T��Z}#��#�L�H���_����+B���