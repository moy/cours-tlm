XlxV37EB    fa00    2252x��=ko۸���+����N�֒��N�8���:I��sq (���%IN����w��$��v�vw�}�4�D����p(�������#�&���;����d��/��l��_�̗�A��A�}`t���[r�0'�n��OHJ��#��g���Ӂ��������w�z�d��_�����!	��	��zg���������s� M�8q�q��#��X#-�x������(���L�-^x�k���Q,��"��g(RQ;��"����޹t��0�|~M��n�JyjG΁H��N�~����#?x<`���v0�Z�{�k���|rD�����3׻M���"<H�o�#��!S�;	�[Ϟ�D��ޱ���xꏿw`���oۻ�5q�����J jYTp
��%��xN�������֎�m�M&΍�9=Ν��_}�p*�#�y2y���s"v�@ó0��x0���o,���k׳A�\{Z�(��τ�sw�L��� �|�H�<�%0�q�p�a˲9��{ю*`���NQg$���{�Ŀ!�"�/"2��H���&��c�O=�6"[ f����j��k��G����8�;��Z���0t� ./�OG#yj羇b � 3�6SP��o��W������_�������k7[S�:��G�:�s�
B����5�oݱe���t*��3�>�;	�3w��S�OǺ�X��e�n��/�#z�
5�C.��vf�껭 �Z��M�bၙ�1�����������K��u�!�b�X������%qí� ���ʱ5�.>	�s@�:�9xC�ä��l�~'�G�Y���������J�����}���" ;���6����5��tَW��w�W���m�l0�J}����S�?:ퟜ\B�T�1X�F�D>iMD�e��?�
���w�Ah�e�B8����|Y��V���`�YG��Q9�zq?>�W���%��;F��(��8:�ގ��bТ�rU<����3F�`8����������DԻ4⶷S�:u����t�e�4j�w�}��,h���"�`��V2	X�i�{�h2d�?����P��}�����_:��Q�>�����Z�ku0p��`T���
I}ά>2%Gːr��
�)4"9�1�>'����}�^򁟽��=*h8Q�XD^���vn�����Q���E�y�F]E"���� �U_�7s�	�?n�X�Y�u�
�#��^���.��d�Tm�ލr$i�T�����4��U4g2˩������b6�艔�"������{�>�q)ћ
�)U�PcUԶ�*�҉��6jӥД�����t�ai� ��)�:\K��`94BB��V�5ǉ��ep��Tiи�K����pp����P;T���q`	��,(O���- ��	���a\L���]���ޠA�# *�����9���]6cj�A!v���d�q�p(ݻ^�^�*����G爀�����=MXS�/���ýu\���hxF���{C\%�T/�C8g:[��~�s����ߠ����[IҌ��9���H06���q�p׽���M֡4P�Q�#C�a�<��<���E@d��=��x��#���������`fܯ�6��όgc]�G�*�X�F�lfx�p�PQ�O������4֖&<���,v�+��<	B�-:�Ⱦ��]���C��Seu���)	S�p������^�p6)eqR�e$]:�o1�>��A� v�:aH 1���Ё6��m��mRH3�[�f)<���U�w��� �p�g!��Ɗ3{>G�ޤ
�E�'���/��m<@�h\X�=f2K�&��H�a*�
�w��	��n"��0����=��M9JY c�#�Uc��h���!����[��3dNr�C��{hIWK�W>n,�:4c�}&U8����E���6nC�{'@G{c�S�P�Y��m
���w~WRԬxcQg�/1�ܝ�?uu:g�:򦏔c�� rv��=u'T@;p� +���@S�� @�~����M� �Ƒ�o�@��:��4�O��찟��-m��uy�����>�z���eztr::�|�\��4m�l�����9V x$�6���Ύ�-���/`F?9c)B�9�W��gh���X�	��u`�3]:�t�n Q��y��8���F�{C>.�N��M�4�?\^dn�>�/����>��dҊr0��Q�N��!f��͘���0�oR���	3�&�.��  I�,��Z*:��~	fF���]�g��)#�W@�Y�c����-#�S@D�m��~�L&�˨0��T�b�իv�P�˥���W�P�P����%%��QN�'D��P�S+%����1r-`�@�u�3_�� �X#���>���' %#
Xm|[�q�n����uP���[�,����+
IƦ�ܹ�����f9��"�	�����e�,����Op�.�D�)A�-;D��N-R�(`��o)i�}��N���h>F�YGwfG�v��N�8:�j��*�c�v��k��:��[;�nV?�gV/+�U5�l1�Y�Ucd��k��������$5�I8*j��pT��'ᨨ�O�QU㟄���k��o֭�=�Ѯ_�{O�)�]A�6�W������~e�_�{�W�����P�^�����󎂪~5W0t��r�a֯�*����\Aa�A�U���\Eѭ_�;��q�Z�U�<�#��N�Zn*�R����ۑ�Z�`د_���-UEW0k�q�	ư���(:���{[U����f����}���l+�խH���®5��W�SU��2�WkX��n	���e�װ*_��V^�?��d�ۨ2��l&����1��� ����xs�h��n��ұl�\�&��Wpt��vn�������W͜�ryP���7!�a�X�T`Ϡ���E������V�I�zƊ�JA� 5��$��&�7e�=�HR:�����PRǊF5�a���\?���M����޳�֎b��ܦBI�v��4�Z$�:g�e�AY�Y�~��$��y(U����d��MY���.Z_ķ5���d(�8�vA��j���Ɣ��sVdh<^?��RY��H�e����#�{b	r�΄��{���5[�!��7��IXnN����c�h�=�P�td��S�<�m�%'�ŋA�D��X�C�ί��
�� ����Z�qUE�记F<AڛdG���CBk�@��4:����?���Α{�=�U�OъFw�Кt�Y�Q�R�=ߨt���F�w�vMG�������I�I&J�JE���`	��n�[��0�&>:�7
�0?[�p��@���!�gb,�:7�#�d�U����.�x�Dx�]��3�w�b��0��8�\�@�A��λ�l~Gѥ��x^S�>'��QjJuCl�-��e>��C3�"�{�W�-�O�M|??�%���'Ԗ�8w��#���U�=�@Uz|���ƼnE>�ě�RKm/=�m�er1��1Y��̿G��
]v~�����_FW\��lo2u�Ii!/:Fvd�G1s�h+Շ�*��:���bF<g��/�w�"��X�sV3˿ǖ~������-h�����eR�����KX��� IjPcKM����-L�M׎��6$��&�t�]�:S�iReL�Z�v�����`�����fy`����GX�����M,���`1�C������Xx�7�i�L�rxD�xT:���1���Gtp]�v�z�"����#-I��vC�U� �4Wh۰�r1e�N�9��jL��'��S'�:)i�
K�i� �wfpCbO��=,�n��E�8��~���0��~xA:ύ獶���3:x����i�++���D�o�mN;8nht���Ʀ�"A&��-�ڮ6�WtT��Q%R�UK�{�s�V�N�H��7g��K�N8"V�6u�~�e�1<�w�%UYb��tܯǝ��v���p;�같lg�ѿ���d�|u'��~N'j_�;�-��iR�~��FR�!s���_]!��X<%U�c���b��/d� dq5�䝥�i�#������O[�ŉ�%Ą�B��lA���8��.I��c.%�8r0���0����kfV 2�L� L�apsU�RR��`�2|i�̗��ҫ��t�U%�*U�̈��nWDۮ��h;+�-��W+���o�愱�Nl5^����M,���J3�*���?�/�Cr��D��{�
�'|9��?�$��E�	^�@s,ʃrpȳ�3��b:���3C�Ǝ&*��篓�;�L��f�W1m����>�$��^~�}>�I�����������.=	�Мo����v�r���y�:`'���)�;g��KO��7e C��������Q&E�����HK��g�X��f@��@m��|G�cK~��w�DB����7��j�3Kb�*�Ͳ����ü�\�t��O�k]�NA�O���o�@~�o/0��\��H�`"؜+����A���Y���7�-���?�-�9�A;ي쥏t�17���1�to��Ya�n�1`�Ē�d#�@�JwpS����͓��;�������� 3�>���;�� [����Cg��?Q��g���p8�3�~�
�������>�/�����v�L��� n�]��Z}���b�\���[���Jk�=��X�8ct/,�ix<��OW�:�� �7~4؂ڌg����Y^�e�~>�����{2�}������i�2�{����}�'�:���"p��L�O�l�T�^s�,��y���7jv2uO�+�6F� ���>����k#�ҥ��dE�F��~����#�AI���hui>z�4��~�nei�}�ݿ�'K�Q2���`�I��d��ń�(����v�iXQʏ��G�$�(�d���4��h��b�w���D�[�'�%}�ѥ�}"������5��>�xU�'�U|���OlU��e|b�1���,L���y���u����O{������Y��,��� ߙff>��L��
�8�Z�eY�Z��:W�'9W�Q�k��o�-�Z{���X��ƭ��j��|]٫U�����X�Q�L��j��/�a����Op�A�;-���8�Z��~�W��|G*ͷ|�VZ�n,�C_��B[?Ʌ���S��v���� ]Ƀ⅍�'x��$W�n5�6Vpy��`g����G��Z2�5��ҩʟd�;Y�mV��撖���Dˍ6���`�ד�b�*jh�`�iV�x����˭�}=1|="�t�'YnS�%TeGh�!�O���6�����4�~55l/o�i��&��mv��+
�b���e���ʐ����JEr�[����bM�3��5����A� ����/��\�v�� n\ܦP����I\��[c`����W�l�Z�/�	Qf���?u7�}?��O�m�Z�����M�����������G�����Е!z.&�^���������Mm�O�|��7��]�Dp��K��5x;��Ij1���cNdP[����.�}�V.�T�'��)|����l���n�7N�oTE({�M���H��:�wGo��r�)%ܘ�Q)�l�7��?�|o
	�4�f��S�ݧM=�_�|?�?�����	%�'��{SMX׶DQEa\t��Q*�g*E���G"���h@��T������9��'#&�^�s���;sr���{�۞!�����	�������?�Wx"l.vl~�y�� ݎ���^�|���س0z�:�� ���aY?� ۔PN���k|�06ݮFA�a-=��S� ���l��ϥ\�/=�X���eEd�c'A��ߚ���g��M2ݕ��O�=s�/����kf�cN^����d��%��Vv�n��F*�����z�L�a�柩�go��Dh򝎧�`�#��	��L��s1z� �b���9�"��Gw��\�R)UIj�"i%9�l�vA��$&ۿV��>�!u�u|��lR�b�W�"��2Y����g�����h\n�Y�6�?vf��O��G�k�%=�Ѣs���3#���nd�8�p ���{Fva������0��u����W����}�P�~l�V:�p	�^�[�.��;'���un����։h,�Ø�7Pe�m�k���Oۇo��`xvd��}|��ŷ��pe�
�y�%��K�9�Qx�|c@%��ߏ�0w�3�<ƞ^�A��n�!\�jv�ٷ�V�:�d�Y��-U�h��v�%}�ܭ�uD�Af�n5��V��r��Z��U����	��W�E9G��7���	1�˟4i��UC|���#��H'[��5�)z-�]]�+*���հY����Ů��N�q�e%Wgu/�ʚ&�⁢}ȼ�/�a$I���e$(�vW0qǊF"~]F��㜜��Hd,Ab#N!�\�H�6Fbc$#��
otx�jj���4�-�����M�%���_ȃ�8��.w#��'GQ)c]-���u9�mփq	-����ķ"��2���;ce��5`w��L�!�e��US��i�N�vZ�J�y�GO�4�W`��?uT��p"4�|'�a����0�"��y�c�6�`m�%Olp��G�húÜz��om�^�WC��^��󪔗���_�~DM��_"]�L���yǂDu�U9�W5wY5I]�z�$�.�����^crz���R�駊GՉ����6���t6!]���,���P���#-y���ڷ�Ji;*��"?~�.ӕN�&{�h6Ѹ,��E�����x��NЙ:S0���\|8�n����0
J���@:�7���7_D�YR%�S=�.�?Z������bnTv17w����5K��Y����*;t�����4�^.y�od��2�#犌����뙻3���ϴS߼I��l�m�t��D$2���&G������=��/�zJ�]�N���q�&����
3f<�7Ԗf�ғ�C��h���:����Z�cX:�D��s�N�"���r�,���,∼�(����.�(�K���u�TgÇ��Jd�<x��:? �p�H�k7�]�c%�M��K't�o��O�5��CR����7�|�_�$��8r�r!L�y�	!o	���gd��S� G} �8Ƕ�`ӂ�@�N�"2�FtgS�م�-�z��0<T����D;��p
�b�%�,'�ʌ�C��N)y��f�Gk��e��2YU��{;p��c�l�5+�	$
@r],|��Nؔ���4-%I�\���g�x�s��
ˤA��1�Qt��X��)��ge�Ѳ]�����e�|�Fe�+�2�H�uU;�X�!JWuj�N�h?�{�ڬ0v�S�X���M.��6��
Ua+8fA=�:�i�����
���kL��.��V����WN���^�Ӣ&4�`P�[%����9��H�R���λ�3cl��h�f���s�yp�(� �d����2��5T&iV��b9�4���%?Xb�v/�X0���l)�նR�r��Q�3��m�ȗ�!AWwB�bm��dx�JB�td��e�'L5����#j�x#+I�Qh������<J!
X& L��:�S�	p!7���g?��J-�n}���_f@�t��M`"4���?-Y
V \\G�s聎�y��N1���(Ix�s-���'� 
�d8^`�7�����<C�P�ɮ�ї�ѾU��"QHw�*pPF�l��p*���ǵ	"а-ˇ�.yN���ev������'3˫9�L��]Q��t�[Q�oH��֝�5�r2-=5L�:�Oi�e��#2)T��f�
)D���� �`�
p�o�y�8��,ה .�6���S�HPfl���"?��gSǻ��O!E���'%#F���������@=7TE��b���N$*3ђ��S�SlY�łJ7=���Q��{�(x&�&b���x�d��gd�+�2W��W��/�ʨn)��=��W�n<SX����ϑ�xQ{�赆 ���	�xPXO�G ���?���z�O�ӷ$4���b}#�6�Օ��U�p�~L����5�^=�Κ�#@��R�el���%�CL�Y1�!�R�DӰA`?6bc�ޭ�Rn�Ύ��#�YWBA�%Le�3�=/+E0��Tn�N%,4�������qܧ��*�ES�t�U���<��I��#%��Me_]%��z��0�sǙ��N���Hs�l[͡�	}����v�ȟ�@�3�|j�����'o�V��l���0��S����A�Ld�f[�mh]��}�j��e��D��T��D��0U�[��Fw0��4RQ��'�5�!n�,�ѧ	�>�����q��ٓ��ޓ����|�1w	㞹�;õ>�ʍ�a�τ-ɼӎ#0v^b9����Q{>��ČZ�J7J���P�Z/o�<��������~�_���]��8�Ɔ%�T���4YP6�v��q�n�72��2�%vA7�u�]��\�>��?h��t���m��o�޻�j.,��[l��#��c��A���90A�LZi��K�����6lo�k����F��!�ǉą�cY�<������y��2���Ǡ��5��]��9�gq�+��q"L�'8?��'��G_�yy���
F!,Y

��*NgzG��C�8�rg��q�T$+��+F�b�5�& �*���a�
�?�2vXlxV37EB    9199    11c1x��]mS۸�ί��Ò��;)�rg�h��eBض�Ύ�$<;�8�����/�,ɖ���Cqt������ ��h�vgh�{S�\���|�;�������m���&�����g�\�g(���O�}o;@����=�'��Ai���5���8F��.���è��h�������b`���kx ����0�����''ck�=�M(�/�y�˽.N�L��	����es"�=x��I��i]�[랮����o����C�շ}�������k�:a�=wf����·�l�ݙ;�w��ww�}�f�����Y�:�Y���;�	����1OF��ط�	�o��>:�u�<�:2�!r\�$#��g�;��}��Y�7֬b��A�;�� ������pF��͗�Wk���-���-��HB>]�e�9��3X�º��0ֿ�:�g2���6��?�m��k-!CC*~�[��y�:�n��2[�_-m��T�Ѱ�����*z��b�������?��$V5�V�h�f��g�]�v��Yٰ�Z����4�ajN����F�D��'{�j��N�D,��݆(60��9�e0��޽3��#�SRއ@:��T��z��.%�Ry���*`I#Z��ƞ#�D���Y(��gQ���\��kjy�:F������������r�`��s��X��G�n��S����X�K��M����z�k;��{ʿe�MT-xxz�\Xh���З��%|9&��e�[�#���5|Yp�D��o����f�/�;.o)�ԈyHD{$��8�up�4JG�
H_��-�m!��hEȤ�����	"S첑�1z���TN)��(k�̔*�����ٸ�!��72?���vܺ��}���s��jA]���=��mJ�8�`�/5lE��BU3'Te(c�6��E&��|I���Q[�MK���Y⹑�RX;����,I:%�W�T�����C;Wd� g3�	8\�� よl(YOE�*2_�������A�5�}@
.�`v���1�j|��pk���ͺ��\/HS��:lI���E\!�6$�W�(�0��^:����rL�Q~�z)57А��!�j�
S� ���(�:K�F��4#^�AVQ��|�Y��L#Fj�|��%m7c{��rˢ%e�(�]�"�9�p�E��U�����<�=�}x�jʋ��W����&i�w���.��k���$n'��D�^��x��f<.�0N2�-���h Y�D�v�f�.q�Y���h?�$�t0`Ј�0��z"�o��طs�����4�zd}����k4}n�M,�S�z�����+ ��Y�N�8&.ON��o��7�ks��-�k��DF.#���?3�C�Z�<�K�K��]��뷉�Q����V�t��0�<��9;��7��U��t'8�p=�hgkУ��:��G���C0��3�����1s��H$�,��=�k+��xVK�b?5�У/V�g��oوfP�����1�;����M֩rv膯c~q#b��}J�d|0�-ѓ��i1w�`3��/|0?r4C| ��P�R����S:h�,�
5��y0�9��1B˕;������$sD�<�&~:����evY91���G�'H,�����?qJpɛr��!���qHG���fb}�p#Dm�_ak�$�&a�$���� N��`���(dʚ��m�sߛ��l`�`�%��� �x�˗J��_f����X"�;��L-��8�)�Q��U�A����c��i��X�?��o�M^��t  �L|�,�h:������!�����ƒ(q�Ý>��뭖�m��i�|#�~�Pg��"+9gYc���b0,n�2��A�P��R� Z^�q���+A�I���<�v+��� ��*���hIf�
����/��i�ͨU� m��4h�v�y:�%���b�i	H��(�!�:i����؎�SM�1������eF&��,*ʢXɏ�������LmE%P�4��������e"F���V������I��2/�3m'lϹ����ur?ԖS�/gZ�[[�Va�v^1�N�,2����0tVX��Zȶ�kV�����C�G����*�c�<a����P����R�Ģ�h�]�����h�=�4%C�)��͒v���Z6�^ͺxn��K!����y>Ӡ��6�Z�;\�K*���=�������h�=Ev�q��ɰP�Z��RY���Gd3tl�9lu��na����"���%4zh��4�"mʒ�F]׻R����Q���ԫ^Vc�FfE%j�I.d��q+<"�r8��En���*L`���r���֩�EX�Mc)�Z��P/�戜��/�#��e�U�Bl�&s�{��j�dd��uEaL��J�ʷ��I8��%IƸe*��u����w2�R���o�۷d�M�qd�N@ݾ�FBqN<��zŏ��ݠ�r���yy����|���ꍻ�q�Y�9k�}8���d��$ϯƗ�[�W��{�Rд�u��j�f���8�����P���-C��9e����H/�δ�%�^~�ܟc۵nt�`�5V>��hb�u��L�5��a�'�
��<n�����3��cs$�C�Qlj�'�XR�pÑ����Aª&<c�%�Ǉ�rM2�gTF!)e0ՁfWg�y 9� ����;$A��`A.|}~���� 1I�_/|�����e��8�Г��A*g`"�����y�n�V�p��GC���p׭�hyAPnǨg�����6�9����5���-(�3�ԕ�*��տ������'b�o��qw2��X���oĢ���!�}~y2���d<�X�����Mt�"" �?�H{i�z��@&,�醧�!&�KU���Z��	�^ď_���	�n2�vi5�]O6RLBlk�f=����*>b٭$@!m�4��A�o�m�/�}kh�^_��e��^Y���S�/�R��W��씻qe,���;ٶ�ɲz�Op+�M;Ĺ���\F�vM��L�5/#���mdT�i�\=�/|s���aJ�bJ��LRg-L��(.�ό�6n�"�etȿׁ[k}�D�<�fh`����h��=# �`����2��)�52��[33����倶�E�-���0�v7C�M�ːP��r��q���OD�j�[1����(��FG��Cm8=,�������tS(�I;:����vB7���v��� j茶Y-�v���>���܂�<U�i4s"��f�9���-ǃ�Ղ��갳�S�Ӭ3��0�P�̶6d��@f����@fYId�C�jﵶ��-�����ͼ�!�l�_)��J�1��\�-)�z�fO'w���3�#�}y�� Ue��t>���ָ���ʀ�u>�;��@x3�4�(�Qp�R��X��T��{��g�k̡U�6�|p~9�jM�^d�cGī��^ٹ�@�_%�.�ͬԍ/#��p�Ny/����P6]�P��pu��L'I1�p��}�@)3�!zΜ�����wi?&>q��?�y+�y��r��r�>,�<l3ǐ���)�j��P�6u]'��D�6��:��71�����;/X.��Bz���F�
u�I�{:�Ͻ��tm�.��E���ܺѿ��M�H"��Ι�/��y|�,"���պҙ���mo�l�U��U�U��ۓ��|���h0�O*�mn}�i���U��Ct��*G�ʪ�ͩ�.D+Y��̡�J��V�%)�
v�<Oy�Y�D����v���N�@��ѡUeu��L��a���f������Fǥ��l�S{��K4�|��O�;4�)�_���<�)�s(�t�	G� ?�3��~t9d>KE:�Yȯ��MG��Ҥ핥U��4i{ei�4U:�([ٖd�H؟0m���D�C��aE��@�<�h9*�/�]O��f��̎�0�d����l�4��b��h�e���B����l��¹�V:'bo�8xKO��'�0�}�UV�U���%�Ǜ!r՘�*W����BȬWǗ��M+�"p�XX^U�>�B�e��T1�e`y�),��`y�(���`�++�{���I@��ZG����J�m|��#׬%ԇp����U��+��f׬����;�e�)$7r��S����WVL����rB	��C�k�Ayk�[�܂e�*�`iK������V�p!O
�Zf���� �	�[D���D���ЮM����1"�(u�����̪��,�G*�-��,�GF�x!O
��-[��-[�.��U[n~jY��e�C5"Q���ûš-U�C��q�U�xo-��+�>/��;H��).�e_{���b����D��\vK��JR!}ҝt���v$[ꆘH��1~ֽS�z[~�-��7���a��
ѭ���L�k��7Q�L��A��ĸ��#�u�M��[�>B�]�ۆ�-�k�Ws>]ģ���ެ���yrY?.��������W}C/�w7�܌;z��mMr2��P��%���BP������o�|���W����b�