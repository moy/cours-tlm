XlxV37EB    34cf     8c4x��Zmo�J�ί�h�)��$m/4�(!��4�r�hue�@��MV���̌_��6/I�������̜�9Ǟf�E�J���t���e�$�{�����
�'*�Z��w��N�PK뜝uZg(�8�O��q��*͗_Pf-�0�e�\ ��O�=������c�y��=�A ���+b��}��ʿ���9�DkX�#� ���j{���]?{�Ƿ���b�¾�hك��گ����&]�|�k+ʕ����[�{��$��<�ldHVv+���	��#�XLIG^��x��G�1��������χ@m��f�Ÿ\�~@��gӽ���xn�3�	wE\�A'�6��"��~�����	:(����L�3�e:��1,{�&��XM܀�݆h�1�XK�����Y��Q�`K�rd���ѧ)�||w3���i)Asl��䑊G���8s��`�(�Lgz��bp%;%�b8o.��8\>�5����~J���&5��e��lR��.�g����!e`�P"�g�ـ�D o��%],)Zx��I8;�͂ 5	閛P@#�xn��x� M@s.�e�{t�X������	ًl�˸��F��i��� ��\Lm,4�4���;�n|z�������OǞ��B�`0�V @��I@-��f�i�����8Ҡ����3�H��\�ۦ�M�/b�N�V������?���Y$&s��^8)Kl�I�J�T��j�ƾ1��ƨ�čq���_���r���ǳ9F��r0|��t�o��P�%U�ꜣ���jC7�w�G��������)D|�=��	�B.X�.iڶ�0J1BܞXLD>ƒPd�1!��Z�z󦪈�z���G
�q�y@H.tC�L�����W�{c�n��V�x�Ay�Q����b�(Y���|���M�~N��k�uG�+t�(�.�s���^�m�sT��%�hB���3�])qV�<t��g�=l��F�~���Ɠ��<�"�P��N����	!�Zg�4�id�Y�/��R�S���આ�J�x
��Bx
\�T8���`��*D���!�x�]8���q�eu�-0]t�"@UȈ�tՌ-�����E�L)�B/TX�ȨP���S"� �(#��}#�����c��յ�"�x1:"��x�=RK^��'�����<V��+��`�0/j�n`n\�|�1�LQ-��ޝ���J
�T�����0��?�xPi1��=$��� #Zd.��g����%�+��k0��"�WBF`�
�6��Z����ݨ���;��Z���3�#\�\/4r{(&{U�H�9{��n�-w�ɦ���<3��"�Na�~ǭ�Fn5�D�L��?%h_@�=�#.fOcG�婩�QQ���T��3�>$<̵2��Lg�o��.��/�Ӧ��A�.a&��ܐڨ�o��ͪ�vU�(%��^���A;yb���C=Z�^%Ry�DB���n��T.����&���!E4w�?�����n�Jc��,�򾲱K2���o�e�@Æ��V�z�c��MP5m� �RP���4����ߑd��kZ]�b�o�{���o�F�_�Fڇ��H{�����F��s���*s��.H���^PVVn2��x��5��-t�#ݖ�'��Rlm�m�T���YJ��)%Um�(E��Q9U���꿶oOԽ��x���!S�m��$���S{ro�lgR�I)��@5x�Q#_*�E�{k����=��C�|���{>tχ���=��C��?�=�C(���{ڮ�Ĥ8��E�'5�|�.�z�~bf��������*�u<�q���\N�9�Ov ����gԳP.���$����]�'$ ��Xϖ�9�a��s@g��J*"�<l��}���ːJt�#9Q�K��"��9&�0 {~��5~����m���(�5#�������[HN���"�*�q�%�k5��)
�$���#�"�©���Bo��D��<V0�̘+���	��	��J�+�T�>G١���Ը �d�l3i9qƮe�F�OlY�Vط��Z0	v��/�K7KF�|a�b�J�7�;J�Ҋd�ԉ�s���2щŔY�\ ��C�����<!���f��C��d��S��S����v�xF���eQH�Z����S6��m+p	q�7������k*f%鋬�3������S�{��TdM�i�B^�:��l