XlxV37EB    1674     61axڽXmo�H��_1J"5��}����ZBT�k��ju:��`u��owM��~���b09 QD�/�>�3ϼ���^��^��~ҁ��{ݘM��Z�����/[���64۝7o:ͷ`��V������5)��:���nB% L<�cW��F8�ߵ��������wO��W0���JuW����1M��`Т�aҀ��"o/WE��TZpx� ��	�,�F�F�f^�c� '��ȓj�M&��
�x���Y����Q�0a*�W��2Fe�Fgk2kޙ���������\�Ʉz�+��`�U:��0�ʁ��H����G6
��T&K%�� fD�J7]��A{�����D��f�#1� ;bRC�"���y*h��4�|S�&o\��;�o-����,Dı6�T���DPnO�.��z����u�P�Q�%p l]ڃZ�T����r�?��ȹ�,C����-�\����Xh�Y;�/U`����_��
*>,��ӂ�n�ϑ#�����[ć,���@�$Tj�����@���M?�H�K�p!N����g�%�y�m�7Cc���"�,�MK�%�PN���B(U�/0r�x���%i��/J�MD(�`*f��͔Gm�/IH#2���͈�b)B�[*ee�o�w���y��o�Rw�^*�b��6y���,$��������~���/�Gq�4=�e��Ta����d�AnW\xl��m��-[�*N*'3�������9f���vJ���g1✣���9��o���~�p���{����^=��g
?�u6i�n���X��6��yMm�W��L�%St���8{����T�=
O6ͺG/|��f�	����φ�V��~�R.��(���,�w�V3��u��j�T�R}VN�"����88��%�f���݀��ӿ���m���a����`���c�S,�n��
?A�Fƻ���V`4D�\�c_Z�<��_���U���'A/T�����3�����(��*.�و�%���ۉb��*�\�z�h68�p�6�4FW�09\;�P��!���ʝ�*Lܔv�YQ��'�4�*툆Ӽp�B'W�%���&rz���zBў*-$��h��g�#bN���&���4
U��>$�Ը�����]�k�a@VP��������z��������/n.��^*�T��B���E� �Wúd�ꉌ������g˭7�
e6��a=��
�E�f�h��p�A�Á��ׅ��Y�X�XZ�ᑅs��aFc�6�M�p��zˣ>=�}
��)��� ����-wS.<x�ǜ�Q_E�*�/��K+U��Q��)Q����\qQXEST͝/7?.ބ�Et}]��\�7�#6�����-���c��=���}`���G�>l�}X�o0��r{�1�CE�e��2��dz�~)�H�VA�	_J	u͐U���	�{�~;Eŉv�:����0����I�^l���~����8��F�B�<_����YK�M���?���%�"��ސ����|m��<����+��7O�plW�Q�����|ѹ���E�.xl�