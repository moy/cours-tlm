XlxV37EB    1d2f     734xڽY[o�J~�W��H�(��C�J	�'Hi��j��b���볻&A:?���bcsM+�_H흙onߌ�Zm�W�VcGݰń4V����>��	k֛��x��|u~�筷o[�w�Xnזu�vT��N		�����N�!�:�M5T�iv��k����J�Z����}JQx�S�]DB>WYWuvE̝0L�=����WA�N�����0�³e���c�X�U�X��U�;!`�x�}B���J25,{Zeh+�1H-��m�R�f�@`C��ΪKf̧l ,5V��T"�2J�R���B1�d4eI�MʥeV1;����f}�#g�0�G Ɛ�'a��l�w��}��
Ő|6*�`B�D�R��W�'�nq|F��
sS]�o���%�M��2��J�B���|`7�C� ��b�Wƈ�8���75a�>�R��� �Y�I#!��K���2�&�Ҷ�'�1Cq�,��_1=�{f������A��ݕ����`���K�D���!R�YٿƤ`���
$�Rĭ��hn����g�
}�f�$�%섴�qjгPh$���+$B!�i�9���~����f�Ȃ*�T�����)d�Y���K����0$7.I��	�,+��]�on�����	�<�H�|�:}��u�Cc�@��p���"k�?8��lh�Hf=�AD�eq� �E4��x���u�l��\EMeE��;�v��c��$"�<�V������k0�	՞?�[���7��Zo��t�n��z�{V�nk�B��#�L�X����Hဤ'_a"L.���wh�=ra�n1�;�VߣY*n�ٔ�����s�f�����|���o�=y~�c��m%'��!'��p�H�zbF���Mke����A.�[U�s���
��8����a������h-�/Q��"��X��#��E�I�˷�g1\'qC��#;M`��?�;I����+�$�q�Z+bf���ִE.��\P�T<����D[��@�����H r��2�a���|�p�.�A��d0�tr[N�i��)���a
{���^PL��&�en4���Z�M�#A�ؘz��3Ű�έՂ��\9�W��$�RTЦ��M#¸������ʩM��2 
���tQ�}��������ߧǻ�ǝSE$�
Y���\T�?�_uc�~�F"�7����q�^T*�ߵs��Ͳ�Ğw#;��v���r�(5�l1�'py�������c���/�7���ҙ����?�����m���ϸ#�tҕ���u�ѸӆIfsg'��*}Ҡ��u��� �_���e���Ft��):/��Fր�itGg:7h��A:z�Fwt��<sغ�5��0�B ��R��*~�a���D�RC-�_p_|���]��`����d.r��""2=(���������0�C��\�"���O
}xA��z�u;q��4�=�صJ��U*"�}��|q3ܓ(Y�{J(�C�3ӿ3�}	O�2R���8];�����)�
1�eu+T<���9���2��H��O=�����5���{�,p�v�<f���uu|����}��\|R {���
A��%'�a^�&�V��:ө-A�`���!Z����S�v>X��J�p�3b�U��]짒{(���Nq�BK ��ͺ����X>&gu�o*>��+�r�����5��)֥�AK~���U%0��>����R%㓂Rmvї�o���v���,)Xe6CtV�;��ƨ�j���AA�GB|M!�>Wsf=�Ջ�?5�Ǎ�uЋX����a�����}��9#*�Z�򑁅��e��?tfnL